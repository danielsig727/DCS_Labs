# INPUT 91
# OUTPUT 79
# NOT 167
# AND 197
# OR 137
# NAND 64
# NOR 92
INPUT(G0)
INPUT(G1)
INPUT(G2)
INPUT(G3)
INPUT(G4)
INPUT(G5)
INPUT(G6)
INPUT(G7)
INPUT(G8)
INPUT(G9)
INPUT(G10)
INPUT(G11)
INPUT(G12)
INPUT(G13)
INPUT(G14)
INPUT(G15)
INPUT(G16)
INPUT(G22)
INPUT(G23)
INPUT(G24)
INPUT(G25)
INPUT(G26)
INPUT(G27)
INPUT(G28)
INPUT(G29)
INPUT(G30)
INPUT(G31)
INPUT(G32)
INPUT(G33)
INPUT(G34)
INPUT(G35)
INPUT(G36)
INPUT(G37)
INPUT(G38)
INPUT(G39)
INPUT(G40)
INPUT(G41)
INPUT(G42)
INPUT(G43)
INPUT(G44)
INPUT(G45)
INPUT(G46)
INPUT(G47)
INPUT(G48)
INPUT(G49)
INPUT(G50)
INPUT(G51)
INPUT(G52)
INPUT(G53)
INPUT(G54)
INPUT(G55)
INPUT(G56)
INPUT(G57)
INPUT(G58)
INPUT(G59)
INPUT(G60)
INPUT(G61)
INPUT(G62)
INPUT(G63)
INPUT(G64)
INPUT(G65)
INPUT(G66)
INPUT(G67)
INPUT(G68)
INPUT(G69)
INPUT(G70)
INPUT(G71)
INPUT(G72)
INPUT(G73)
INPUT(G74)
INPUT(G75)
INPUT(G76)
INPUT(G77)
INPUT(G78)
INPUT(G79)
INPUT(G80)
INPUT(G81)
INPUT(G82)
INPUT(G83)
INPUT(G84)
INPUT(G85)
INPUT(G86)
INPUT(G87)
INPUT(G88)
INPUT(G89)
INPUT(G90)
INPUT(G91)
INPUT(G92)
INPUT(G93)
INPUT(G94)
INPUT(G95)
OUTPUT(G726)
OUTPUT(G729)
OUTPUT(G702)
OUTPUT(G727)
OUTPUT(G701BF)
OUTPUT(G332BF)
OUTPUT(G328BF)
OUTPUT(G109)
OUTPUT(G113)
OUTPUT(G118)
OUTPUT(G125)
OUTPUT(G129)
OUTPUT(G140)
OUTPUT(G144)
OUTPUT(G149)
OUTPUT(G154)
OUTPUT(G159)
OUTPUT(G166)
OUTPUT(G175)
OUTPUT(G189)
OUTPUT(G193)
OUTPUT(G198)
OUTPUT(G208)
OUTPUT(G214)
OUTPUT(G218)
OUTPUT(G237)
OUTPUT(G242)
OUTPUT(G247)
OUTPUT(G252)
OUTPUT(G260)
OUTPUT(G303)
OUTPUT(G309)
OUTPUT(G315)
OUTPUT(G321)
OUTPUT(G360)
OUTPUT(G365)
OUTPUT(G373)
OUTPUT(G379)
OUTPUT(G384)
OUTPUT(G392)
OUTPUT(G397)
OUTPUT(G405)
OUTPUT(G408)
OUTPUT(G416)
OUTPUT(G424)
OUTPUT(G427)
OUTPUT(G438)
OUTPUT(G441)
OUTPUT(G447)
OUTPUT(G451)
OUTPUT(G459)
OUTPUT(G464)
OUTPUT(G469)
OUTPUT(G477)
OUTPUT(G494)
OUTPUT(G498)
OUTPUT(G503)
OUTPUT(G526)
OUTPUT(G531)
OUTPUT(G536)
OUTPUT(G541)
OUTPUT(G548)
OUTPUT(G565)
OUTPUT(G569)
OUTPUT(G573)
OUTPUT(G577)
OUTPUT(G590)
OUTPUT(G608)
OUTPUT(G613)
OUTPUT(G657)
OUTPUT(G663)
OUTPUT(G669)
OUTPUT(G675)
OUTPUT(G682)
OUTPUT(G687)
OUTPUT(G693)
OUTPUT(G705)
OUTPUT(G707)
OUTPUT(G713)
G712(43) = NOT(G14)
G111(3) = NOT(G24)
G127(3) = NOT(G27)
G142(3) = NOT(G29)
G176(1) = NOT(G35)
G178(4) = NOT(G34)
G180(6) = NOT(G92)
G191(3) = NOT(G36)
G204(1) = NOT(G38)
G210(3) = NOT(G39)
G216(3) = NOT(G40)
G348(9) = NOT(G91)
G645(28) = NOT(G90)
G445(1) = NOT(G65)
G449(1) = NOT(G66)
G511(7) = NOT(G63)
G614(1) = NOT(G64)
I1162(1) = NOT(G13)
G661(2) = NOT(G94)
I1183(1) = NOT(G11)
I1203(1) = NOT(G10)
G701(2) = NOT(G15)
I1227(1) = NOT(G6)
I1230(1) = NOT(G7)
I1233(1) = NOT(G8)
I1236(1) = NOT(G9)
I1239(1) = NOT(G12)
I1242(1) = NOT(G0)
I1245(1) = NOT(G1)
I1248(1) = NOT(G2)
I1251(1) = NOT(G3)
I1254(1) = NOT(G4)
I1257(1) = NOT(G5)
I1260(1) = NOT(G93)
I1264(1) = NOT(G16)
I1267(1) = NOT(G95)
G300(1) = OR(G50, G49, G48, G47)
G301(2) = NAND(G50, G49, G48, G47)
G518(1) = OR(G71, G67)
G519(1) = OR(G72, G68)
G520(1) = OR(G73, G69)
G487(2) = NOR(G71, G72, G73)
G583(1) = OR(G79, G74)
G584(1) = OR(G80, G75)
G585(1) = OR(G81, G76)
G586(1) = OR(G82, G77)
G561(2) = NOR(G79, G80, G81, G82)
G514(1) = NAND(G71, G67)
G515(1) = NAND(G72, G68)
G516(1) = NAND(G73, G69)
G578(1) = NAND(G79, G74)
G579(1) = NAND(G80, G75)
G580(1) = NAND(G81, G76)
G581(1) = NAND(G82, G77)
G726(1) = NOT(I1260)
G729(1) = NOT(I1267)
G108(1) = NOT(G712)
G112(1) = NOT(G712)
G117(1) = NOT(G712)
G124(1) = NOT(G712)
G128(1) = NOT(G712)
G139(1) = NOT(G712)
G143(1) = NOT(G712)
G148(1) = NOT(G712)
G153(1) = NOT(G712)
G158(1) = NOT(G712)
G165(1) = NOT(G712)
G174(1) = NOT(G712)
G179(1) = NOT(G180)
G188(1) = NOT(G712)
G192(1) = NOT(G712)
G197(1) = NOT(G712)
G207(1) = NOT(G712)
G213(1) = NOT(G712)
G217(1) = NOT(G712)
G302(1) = NOT(G712)
G308(1) = NOT(G712)
G314(1) = NOT(G712)
G320(1) = NOT(G712)
G343(1) = NOT(G348)
G347(1) = NOT(G348)
G351(1) = NOT(G645)
G407(1) = NOT(G712)
G426(1) = NOT(G712)
G437(1) = NOT(G712)
G440(1) = NOT(G712)
G446(1) = NOT(G712)
G450(1) = NOT(G712)
G486(1) = NOT(G712)
G504(1) = NOT(G511)
G507(1) = NOT(G511)
G510(1) = NOT(G511)
G617(1) = NOT(G645)
G620(1) = NOT(G645)
G623(1) = NOT(G645)
G626(1) = NOT(G645)
G629(1) = NOT(G645)
G632(1) = NOT(G645)
G635(1) = NOT(G645)
G638(1) = NOT(G645)
G641(1) = NOT(G645)
G644(1) = NOT(G645)
G656(1) = NOT(G712)
G659(2) = NOT(I1162)
G662(1) = NOT(G712)
G678(9) = NOT(I1183)
G668(1) = NOT(G712)
G674(1) = NOT(G712)
G696(7) = NOT(I1203)
I1211(1) = NOT(G701)
G704(1) = NOT(G712)
G706(1) = NOT(G712)
G711(1) = NOT(G712)
G714(4) = NOT(G701)
G715(2) = NOT(I1227)
G716(2) = NOT(I1230)
G717(2) = NOT(I1233)
G718(2) = NOT(I1236)
G719(1) = NOT(I1239)
G720(2) = NOT(I1242)
G721(2) = NOT(I1245)
G722(2) = NOT(I1248)
G723(2) = NOT(I1251)
G724(2) = NOT(I1254)
G725(2) = NOT(I1257)
G728(1) = NOT(I1264)
G181(1) = OR(G178, G180)
G349(1) = OR(G62, G348)
G621(1) = OR(G614, G645)
G521(1) = OR(G487, G70)
G587(1) = OR(G561, G78)
G482(1) = NAND(G514, G518)
G483(1) = NAND(G515, G519)
G484(1) = NAND(G516, G520)
G517(1) = NAND(G487, G70)
G556(1) = NAND(G578, G583)
G557(1) = NAND(G579, G584)
G558(1) = NAND(G580, G585)
G559(1) = NAND(G581, G586)
G582(1) = NAND(G561, G78)
G701BF(1) = NOT(I1211)
G175(1) = AND(G176, G174)
G657(1) = AND(G659, G656)
G658(2) = NOT(G659)
G665(1) = NOT(G678)
G671(1) = NOT(G678)
G677(1) = NOT(G678)
G685(1) = NOT(G696)
G689(1) = NOT(G696)
G695(1) = NOT(G696)
G631(1) = OR(G720, G629)
G634(1) = OR(G721, G632)
G637(1) = OR(G722, G635)
G640(1) = OR(G723, G638)
G643(1) = OR(G724, G641)
G182(1) = OR(G35, G179)
G625(1) = OR(G716, G623)
G350(1) = OR(G59, G347)
G353(1) = OR(G35, G351)
G505(1) = OR(G723, G511)
G506(1) = OR(G720, G504)
G508(1) = OR(G724, G511)
G509(1) = OR(G721, G507)
G512(1) = OR(G725, G511)
G513(1) = OR(G722, G510)
G628(1) = OR(G718, G626)
G622(1) = OR(G717, G620)
G647(1) = OR(G725, G644)
G619(1) = OR(G715, G617)
G666(1) = OR(G87, G678)
G672(1) = OR(G88, G678)
G679(1) = OR(G89, G678)
G684(1) = OR(G645, G696)
G690(1) = OR(G348, G696)
G697(1) = OR(G180, G696)
G709(1) = AND(G678, G89)
G333(1) = OR(G300, G714)
G334(1) = OR(G301, G714)
G554(1) = NAND(G556, G557, G558)
G485(1) = NAND(G517, G521)
G560(1) = NAND(G582, G587)
G710(1) = NOR(G678, G94)
G601(2) = AND(G621, G622)
G616(2) = NAND(G482, G483, G484, G485)
G185(1) = AND(G181, G182)
G331(2) = NAND(G333, G22)
G346(1) = AND(G349, G350)
G488(1) = AND(G505, G506)
G489(1) = AND(G508, G509)
G490(1) = AND(G512, G513)
G667(1) = OR(G661, G665)
G673(1) = OR(G87, G671)
G680(1) = OR(G88, G677)
G683(1) = AND(G684, G685)
G691(1) = OR(G645, G689)
G698(1) = OR(G348, G695)
G708(1) = NOR(G709, G710)
G555(1) = NAND(G559, G560)
G699(3) = OR(G658, G712)
G660(3) = NOR(G658, G86)
G707(1) = AND(G708, G706)
G332(2) = NAND(G334, G331)
G476(9) = NAND(G486, G616)
G600(1) = NOT(G601)
G615(5) = NOT(G616)
G329(1) = AND(G331, G714)
G352(1) = OR(G346, G645)
G524(3) = OR(G554, G555)
G664(1) = AND(G666, G667)
G670(1) = AND(G672, G673)
G676(1) = AND(G679, G680)
G688(1) = AND(G690, G691)
G694(1) = AND(G697, G698)
G602(1) = OR(G85, G601)
G681(1) = NOR(G683, G660)
G727(1) = AND(G476, G645)
G663(1) = AND(G664, G662)
G669(1) = AND(G670, G668)
G675(1) = AND(G676, G674)
G682(1) = OR(G681, G699)
I1(1) = NOT(G332)
G456(2) = OR(G83, G524)
G458(1) = NOT(G476)
G463(1) = NOT(G476)
G468(1) = NOT(G476)
G475(1) = NOT(G476)
G624(1) = OR(G476, G645)
G330(1) = AND(G332, G714)
G436(1) = AND(G352, G353)
G443(1) = AND(G615, G511)
G448(1) = OR(G615, G65)
G453(1) = AND(G615, G445)
G627(1) = OR(G476, G645)
G654(1) = AND(G90, G476)
G655(1) = AND(G91, G476)
G603(1) = OR(G600, G84)
G686(1) = NOR(G688, G660)
G692(1) = NOR(G694, G660)
G444(1) = NOR(G615, G64)
G454(1) = NOR(G615, G66)
G332BF(1) = NOT(I1)
G447(1) = AND(G448, G446)
G687(1) = OR(G686, G699)
G693(1) = OR(G692, G699)
G259(5) = AND(G624, G625)
G455(1) = NOT(G456)
G500(6) = OR(G654, G712)
G589(6) = AND(G627, G628)
G610(12) = OR(G655, G712)
G597(2) = NAND(G602, G603)
G442(1) = NOR(G443, G444)
G452(1) = NOR(G453, G454)
G646(1) = OR(G456, G645)
G327(1) = NOR(G330, G23)
G441(1) = AND(G442, G440)
G451(1) = AND(G452, G450)
G328(2) = NOR(G329, G327)
G236(1) = NOT(G259)
G241(1) = NOT(G259)
G246(1) = NOT(G259)
G251(1) = NOT(G259)
G258(1) = NOT(G259)
G491(1) = NOT(G500)
G495(1) = NOT(G500)
G499(1) = NOT(G500)
G525(1) = NOT(G589)
G530(1) = NOT(G589)
G535(1) = NOT(G589)
G540(1) = NOT(G589)
G547(1) = NOT(G589)
G562(1) = NOT(G610)
G566(1) = NOT(G610)
G570(1) = NOT(G610)
G574(1) = NOT(G610)
G588(1) = NOT(G589)
G596(5) = NOT(G597)
G605(1) = NOT(G610)
G609(1) = NOT(G610)
G457(2) = AND(G455, G449, G728)
G492(1) = OR(G71, G500)
G496(1) = OR(G72, G500)
G501(1) = OR(G73, G500)
G563(1) = OR(G79, G610)
G567(1) = OR(G80, G610)
G571(1) = OR(G81, G610)
G575(1) = OR(G82, G610)
G606(1) = OR(G84, G610)
G611(1) = OR(G85, G610)
G648(1) = AND(G646, G647)
I12(1) = NOT(G328)
G355(6) = OR(G457, G645)
G299(3) = NOR(G301, G328)
G493(1) = OR(G488, G491)
G497(1) = OR(G489, G495)
G502(1) = OR(G490, G499)
G564(1) = OR(G715, G562)
G568(1) = OR(G716, G566)
G572(1) = OR(G717, G570)
G576(1) = OR(G718, G574)
G607(1) = OR(G696, G605)
G612(1) = OR(G678, G609)
G618(1) = OR(G457, G645)
G96(1) = NAND(G74, G596)
G97(1) = NAND(G75, G596)
G98(1) = NAND(G76, G596)
G99(1) = NAND(G77, G596)
G100(1) = NAND(G78, G596)
G328BF(1) = NOT(I12)
G494(1) = AND(G492, G493)
G498(1) = AND(G496, G497)
G503(1) = AND(G501, G502)
G565(1) = AND(G563, G564)
G569(1) = AND(G567, G568)
G573(1) = AND(G571, G572)
G577(1) = AND(G575, G576)
G608(1) = AND(G606, G607)
G613(1) = AND(G611, G612)
G336(1) = NOT(G355)
G339(1) = NOT(G355)
G354(1) = NOT(G355)
G630(1) = OR(G96, G645)
G633(1) = OR(G97, G645)
G636(1) = OR(G98, G645)
G639(1) = OR(G99, G645)
G642(1) = OR(G100, G645)
G240(1) = AND(G299, G42)
G262(3) = AND(G299, G42)
G340(1) = OR(G38, G355)
G649(2) = AND(G618, G619)
G239(1) = NOR(G299, G42)
G101(3) = AND(G630, G631)
G102(3) = AND(G633, G634)
G103(3) = AND(G636, G637)
G104(3) = AND(G639, G640)
G105(3) = AND(G642, G643)
G238(1) = NOR(G239, G240)
G245(1) = AND(G262, G43)
G263(3) = AND(G262, G43)
G341(1) = OR(G185, G339)
G234(1) = NAND(G649, G436)
G244(1) = NOR(G262, G43)
G237(1) = AND(G238, G236)
G243(1) = NOR(G244, G245)
G250(1) = AND(G263, G44)
G264(3) = AND(G263, G44)
G275(1) = OR(G101, G42)
G276(1) = OR(G102, G43)
G278(1) = OR(G103, G44)
G280(1) = OR(G104, G45)
G435(5) = AND(G340, G341)
G282(1) = OR(G105, G46)
G291(1) = OR(G42, G101)
G292(1) = OR(G43, G102)
G293(1) = OR(G44, G103)
G294(1) = OR(G45, G104)
G295(1) = OR(G46, G105)
G286(1) = NAND(G42, G101)
G287(1) = NAND(G43, G102)
G288(1) = NAND(G44, G103)
G284(1) = NAND(G45, G104)
G285(1) = NAND(G46, G105)
G249(1) = NOR(G263, G44)
G242(1) = AND(G243, G241)
G593(2) = NOR(G435, G524)
G248(1) = NOR(G249, G250)
G255(1) = AND(G264, G45)
G265(2) = AND(G264, G45)
G266(2) = NAND(G286, G291)
G439(1) = OR(G435, G63)
G267(2) = NAND(G287, G292)
G268(2) = NAND(G288, G293)
G269(2) = NAND(G284, G294)
G270(2) = NAND(G285, G295)
G231(1) = NAND(G435, G648)
G598(1) = NAND(G435, G83)
G254(1) = NOR(G264, G45)
G247(1) = AND(G248, G246)
G438(1) = AND(G439, G437)
G595(1) = NOT(G593)
G253(1) = NOR(G254, G255)
G261(1) = AND(G265, G46)
G271(1) = AND(G275, G266)
G594(1) = OR(G83, G593)
G599(1) = NOR(G598, G597)
G289(1) = NOR(G270, G269, G268)
G290(1) = NOR(G267, G266)
G257(1) = NOR(G265, G46)
G252(1) = AND(G253, G251)
G713(1) = AND(G599, G711)
G297(2) = NAND(G289, G290)
G256(1) = NOR(G257, G261)
G277(1) = OR(G267, G271)
G592(1) = AND(G594, G595)
G260(1) = AND(G256, G258)
G296(1) = NOT(G297)
G272(1) = AND(G276, G277)
G279(1) = OR(G268, G272)
G273(1) = AND(G278, G279)
G281(1) = OR(G269, G273)
G274(1) = AND(G280, G281)
G283(1) = OR(G270, G274)
G700(5) = NAND(G282, G283)
G133(3) = AND(G700, G111)
G110(1) = OR(G700, G111)
G107(1) = NAND(G700, G111)
G298(1) = NAND(G297, G700)
G106(1) = NAND(G107, G110)
G116(1) = AND(G133, G25)
G134(3) = AND(G133, G25)
G232(1) = NAND(G296, G298, G435)
G115(1) = NOR(G133, G25)
G109(1) = AND(G106, G108)
G114(1) = NOR(G115, G116)
G121(1) = AND(G134, G26)
G135(3) = AND(G134, G26)
G233(1) = NAND(G700, G232, G231)
G120(1) = NOR(G134, G26)
G113(1) = AND(G114, G112)
G119(1) = NOR(G120, G121)
G136(3) = AND(G135, G127)
G126(1) = OR(G135, G127)
G235(1) = OR(G649, G233)
G123(1) = NAND(G135, G127)
G118(1) = AND(G119, G117)
G122(1) = NAND(G123, G126)
G132(1) = AND(G136, G28)
G226(2) = AND(G136, G28)
G230(1) = NAND(G234, G235)
G131(1) = NOR(G136, G28)
G125(1) = AND(G122, G124)
G705(1) = AND(G230, G704)
G130(1) = NOR(G131, G132)
G177(3) = OR(G180, G226)
G650(1) = AND(G226, G661)
G129(1) = AND(G130, G128)
G168(3) = AND(G177, G142)
G141(1) = OR(G177, G142)
G138(1) = NAND(G177, G142)
G137(1) = NAND(G138, G141)
G147(1) = AND(G168, G30)
G169(3) = AND(G168, G30)
G146(1) = NOR(G168, G30)
G140(1) = AND(G137, G139)
G145(1) = NOR(G146, G147)
G152(1) = AND(G169, G31)
G170(3) = AND(G169, G31)
G151(1) = NOR(G169, G31)
G144(1) = AND(G145, G143)
G150(1) = NOR(G151, G152)
G157(1) = AND(G170, G32)
G171(3) = AND(G170, G32)
G156(1) = NOR(G170, G32)
G149(1) = AND(G150, G148)
G155(1) = NOR(G156, G157)
G162(1) = AND(G171, G33)
G172(4) = AND(G171, G33)
G161(1) = NOR(G171, G33)
G154(1) = AND(G155, G153)
G160(1) = NOR(G161, G162)
G173(1) = AND(G172, G34)
G227(2) = AND(G172, G178)
G167(1) = OR(G172, G178)
G164(1) = NAND(G172, G178)
G159(1) = AND(G160, G158)
G163(1) = NAND(G164, G167)
G183(8) = OR(G180, G227)
G651(1) = AND(G227, G87)
G184(1) = OR(G180, G173)
G166(1) = AND(G163, G165)
G222(3) = AND(G183, G210)
G338(1) = OR(G183, G336)
G377(2) = AND(G183, G54, G56)
G382(1) = AND(G183, G54)
G394(3) = AND(G183, G54)
G357(1) = OR(G184, G354)
G209(1) = OR(G183, G210)
G206(1) = NAND(G183, G210)
G381(1) = NOR(G183, G54)
G324(8) = OR(G377, G348)
G391(3) = OR(G712, G377)
G205(1) = NAND(G206, G209)
G223(3) = AND(G222, G216)
G380(1) = NOR(G381, G382)
G387(1) = AND(G394, G55)
G395(2) = AND(G394, G55)
G215(1) = OR(G222, G216)
G212(1) = NAND(G222, G216)
G386(1) = NOR(G394, G55)
G208(1) = AND(G205, G207)
G305(1) = NOT(G324)
G311(1) = NOT(G324)
G317(1) = NOT(G324)
G323(1) = NOT(G324)
G378(1) = NOT(G391)
G383(1) = NOT(G391)
G390(1) = NOT(G391)
G211(1) = NAND(G212, G215)
G221(1) = AND(G223, G41)
G228(2) = AND(G223, G41)
G306(1) = OR(G47, G324)
G312(1) = OR(G48, G324)
G318(1) = OR(G49, G324)
G325(1) = OR(G50, G324)
G385(1) = NOR(G386, G387)
G393(1) = AND(G395, G56)
G220(1) = NOR(G223, G41)
G389(1) = NOR(G395, G56)
G214(1) = AND(G211, G213)
G379(1) = AND(G380, G378)
G384(1) = AND(G385, G383)
G522(3) = OR(G348, G228)
G219(1) = NOR(G220, G221)
G307(1) = OR(G719, G305)
G313(1) = OR(G47, G311)
G319(1) = OR(G48, G317)
G326(1) = OR(G49, G323)
G388(1) = NOR(G389, G393)
G652(1) = AND(G228, G88)
G218(1) = AND(G219, G217)
G392(1) = AND(G388, G390)
G202(3) = AND(G522, G191)
G304(1) = AND(G306, G307)
G310(1) = AND(G312, G313)
G316(1) = AND(G318, G319)
G322(1) = AND(G325, G326)
G190(1) = OR(G522, G191)
G187(1) = NAND(G522, G191)
G303(1) = AND(G304, G302)
G309(1) = AND(G310, G308)
G315(1) = AND(G316, G314)
G321(1) = AND(G322, G320)
G186(1) = NAND(G187, G190)
G196(1) = AND(G202, G37)
G203(4) = AND(G202, G37)
G195(1) = NOR(G202, G37)
G189(1) = AND(G186, G188)
G194(1) = NOR(G195, G196)
G201(1) = AND(G203, G38)
G224(1) = AND(G203, G38)
G225(1) = AND(G204, G203)
G200(1) = NOR(G203, G38)
G193(1) = AND(G194, G192)
G199(1) = NOR(G200, G201)
G337(1) = OR(G224, G355)
G356(1) = OR(G225, G355)
G198(1) = AND(G199, G197)
G335(4) = AND(G337, G338)
G433(1) = AND(G356, G357)
G400(1) = AND(G335, G57)
G412(2) = AND(G335, G57)
G413(4) = AND(G335, G58)
G604(4) = AND(G433, G524)
G399(1) = NOR(G335, G57)
G404(2) = OR(G712, G413)
G398(1) = NOR(G399, G400)
G406(1) = AND(G412, G58)
G411(1) = AND(G413, G59)
G414(2) = AND(G413, G59)
G529(1) = AND(G604, G74)
G550(3) = AND(G604, G74)
G591(1) = OR(G592, G604)
G402(1) = NOR(G412, G58)
G410(1) = NOR(G413, G59)
G528(1) = NOR(G604, G74)
G590(1) = AND(G591, G588)
G396(1) = NOT(G404)
G403(1) = NOT(G404)
G345(1) = OR(G414, G343)
G523(4) = OR(G348, G414)
G401(1) = NOR(G402, G406)
G409(1) = NOR(G410, G411)
G527(1) = NOR(G528, G529)
G534(1) = AND(G550, G75)
G551(3) = AND(G550, G75)
G533(1) = NOR(G550, G75)
G397(1) = AND(G398, G396)
G405(1) = AND(G401, G403)
G408(1) = AND(G409, G407)
G526(1) = AND(G527, G525)
G358(5) = AND(G523, G53)
G363(1) = AND(G523, G51)
G375(3) = AND(G523, G51)
G532(1) = NOR(G533, G534)
G539(1) = AND(G551, G76)
G552(3) = AND(G551, G76)
G362(1) = NOR(G523, G51)
G538(1) = NOR(G551, G76)
G531(1) = AND(G532, G530)
G372(3) = OR(G712, G358)
G432(4) = AND(G358, G61)
G361(1) = NOR(G362, G363)
G368(1) = AND(G375, G52)
G376(2) = AND(G375, G52)
G419(1) = AND(G358, G60)
G431(2) = AND(G358, G60)
G537(1) = NOR(G538, G539)
G544(1) = AND(G552, G77)
G553(2) = AND(G552, G77)
G367(1) = NOR(G375, G52)
G418(1) = NOR(G358, G60)
G543(1) = NOR(G552, G77)
G536(1) = AND(G537, G535)
G359(1) = NOT(G372)
G364(1) = NOT(G372)
G371(1) = NOT(G372)
G423(2) = OR(G712, G432)
G229(2) = AND(G432, G62)
G366(1) = NOR(G367, G368)
G374(1) = AND(G376, G53)
G417(1) = NOR(G418, G419)
G425(1) = AND(G431, G61)
G430(1) = AND(G432, G62)
G542(1) = NOR(G543, G544)
G549(1) = AND(G553, G78)
G370(1) = NOR(G376, G53)
G421(1) = NOR(G431, G61)
G429(1) = NOR(G432, G62)
G546(1) = NOR(G553, G78)
G360(1) = AND(G361, G359)
G365(1) = AND(G366, G364)
G541(1) = AND(G542, G540)
G415(1) = NOT(G423)
G422(1) = NOT(G423)
G344(1) = OR(G229, G348)
G369(1) = NOR(G370, G374)
G420(1) = NOR(G421, G425)
G428(1) = NOR(G429, G430)
G545(1) = NOR(G546, G549)
G653(1) = AND(G229, G89)
G373(1) = AND(G369, G371)
G416(1) = AND(G417, G415)
G424(1) = AND(G420, G422)
G427(1) = AND(G428, G426)
G548(1) = AND(G545, G547)
G342(1) = AND(G344, G345)
G703(1) = NOR(G650, G651, G652, G653)
G702(1) = AND(G703, G645)
G434(3) = OR(G342, G645)
G462(1) = AND(G434, G67)
G479(3) = AND(G434, G67)
G461(1) = NOR(G434, G67)
G460(1) = NOR(G461, G462)
G467(1) = AND(G479, G68)
G480(3) = AND(G479, G68)
G466(1) = NOR(G479, G68)
G459(1) = AND(G460, G458)
G465(1) = NOR(G466, G467)
G472(1) = AND(G480, G69)
G481(2) = AND(G480, G69)
G471(1) = NOR(G480, G69)
G464(1) = AND(G465, G463)
G470(1) = NOR(G471, G472)
G478(1) = AND(G481, G70)
G474(1) = NOR(G481, G70)
G469(1) = AND(G470, G468)
G473(1) = NOR(G474, G478)
G477(1) = AND(G473, G475)
