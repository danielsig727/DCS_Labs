# INPUT 1464
# OUTPUT 1730
# NOT 7805
# AND 5516
# OR 2621
# NAND 2126
# NOR 1185
INPUT(g35)
INPUT(g36)
INPUT(g6744)
INPUT(g6745)
INPUT(g6746)
INPUT(g6747)
INPUT(g6748)
INPUT(g6749)
INPUT(g6750)
INPUT(g6751)
INPUT(g6752)
INPUT(g6753)
INPUT(g84)
INPUT(g120)
INPUT(g5)
INPUT(g113)
INPUT(g126)
INPUT(g99)
INPUT(g53)
INPUT(g116)
INPUT(g92)
INPUT(g56)
INPUT(g91)
INPUT(g44)
INPUT(g57)
INPUT(g100)
INPUT(g54)
INPUT(g124)
INPUT(g125)
INPUT(g114)
INPUT(g134)
INPUT(g72)
INPUT(g115)
INPUT(g135)
INPUT(g90)
INPUT(g127)
INPUT(g64)
INPUT(g73)
INPUT(g5057)
INPUT(g2771)
INPUT(g1882)
INPUT(g6462)
INPUT(g2299)
INPUT(g4040)
INPUT(g2547)
INPUT(g559)
INPUT(g3017)
INPUT(g3243)
INPUT(g452)
INPUT(g464)
INPUT(g3542)
INPUT(g5232)
INPUT(g5813)
INPUT(g2907)
INPUT(g1744)
INPUT(g5909)
INPUT(g1802)
INPUT(g3554)
INPUT(g6219)
INPUT(g807)
INPUT(g6031)
INPUT(g847)
INPUT(g976)
INPUT(g4172)
INPUT(g4372)
INPUT(g3512)
INPUT(g749)
INPUT(g3490)
INPUT(g6005)
INPUT(g4235)
INPUT(g1600)
INPUT(g1714)
INPUT(g3649)
INPUT(g3155)
INPUT(g3355)
INPUT(g2236)
INPUT(g4555)
INPUT(g3698)
INPUT(g6073)
INPUT(g1736)
INPUT(g1968)
INPUT(g4621)
INPUT(g5607)
INPUT(g2657)
INPUT(g5659)
INPUT(g490)
INPUT(g311)
INPUT(g6069)
INPUT(g772)
INPUT(g5587)
INPUT(g6177)
INPUT(g6377)
INPUT(g3167)
INPUT(g5615)
INPUT(g4567)
INPUT(g3057)
INPUT(g3457)
INPUT(g6287)
INPUT(g1500)
INPUT(g2563)
INPUT(g4776)
INPUT(g4593)
INPUT(g6199)
INPUT(g2295)
INPUT(g1384)
INPUT(g1339)
INPUT(g5180)
INPUT(g2844)
INPUT(g1024)
INPUT(g5591)
INPUT(g3598)
INPUT(g4264)
INPUT(g767)
INPUT(g5853)
INPUT(g3321)
INPUT(g2089)
INPUT(g4933)
INPUT(g4521)
INPUT(g5507)
INPUT(g3625)
INPUT(g6291)
INPUT(g294)
INPUT(g5559)
INPUT(g5794)
INPUT(g6144)
INPUT(g3813)
INPUT(g562)
INPUT(g608)
INPUT(g1205)
INPUT(g3909)
INPUT(g6259)
INPUT(g5905)
INPUT(g921)
INPUT(g2955)
INPUT(g203)
INPUT(g6088)
INPUT(g1099)
INPUT(g4878)
INPUT(g5204)
INPUT(g5630)
INPUT(g3606)
INPUT(g1926)
INPUT(g6215)
INPUT(g3586)
INPUT(g291)
INPUT(g4674)
INPUT(g3570)
INPUT(g640)
INPUT(g5969)
INPUT(g1862)
INPUT(g676)
INPUT(g843)
INPUT(g4132)
INPUT(g4332)
INPUT(g4153)
INPUT(g5666)
INPUT(g6336)
INPUT(g622)
INPUT(g3506)
INPUT(g4558)
INPUT(g6065)
INPUT(g6322)
INPUT(g3111)
INPUT(g117)
INPUT(g2837)
INPUT(g939)
INPUT(g278)
INPUT(g4492)
INPUT(g4864)
INPUT(g1036)
INPUT(g128)
INPUT(g1178)
INPUT(g3239)
INPUT(g718)
INPUT(g6195)
INPUT(g1135)
INPUT(g6137)
INPUT(g6395)
INPUT(g3380)
INPUT(g5343)
INPUT(g554)
INPUT(g496)
INPUT(g3853)
INPUT(g5134)
INPUT(g1422)
INPUT(g3794)
INPUT(g2485)
INPUT(g925)
INPUT(g48)
INPUT(g5555)
INPUT(g878)
INPUT(g1798)
INPUT(g4076)
INPUT(g2941)
INPUT(g3905)
INPUT(g763)
INPUT(g6255)
INPUT(g4375)
INPUT(g4871)
INPUT(g4722)
INPUT(g590)
INPUT(g6692)
INPUT(g1632)
INPUT(g5313)
INPUT(g3100)
INPUT(g1495)
INPUT(g6497)
INPUT(g1437)
INPUT(g6154)
INPUT(g1579)
INPUT(g5567)
INPUT(g1752)
INPUT(g1917)
INPUT(g744)
INPUT(g3040)
INPUT(g4737)
INPUT(g4809)
INPUT(g6267)
INPUT(g3440)
INPUT(g3969)
INPUT(g1442)
INPUT(g5965)
INPUT(g4477)
INPUT(g1233)
INPUT(g4643)
INPUT(g5264)
INPUT(g6329)
INPUT(g2610)
INPUT(g5160)
INPUT(g5360)
INPUT(g5933)
INPUT(g1454)
INPUT(g753)
INPUT(g1296)
INPUT(g3151)
INPUT(g2980)
INPUT(g6727)
INPUT(g3530)
INPUT(g4742)
INPUT(g4104)
INPUT(g1532)
INPUT(g4304)
INPUT(g2177)
INPUT(g3010)
INPUT(g52)
INPUT(g4754)
INPUT(g1189)
INPUT(g2287)
INPUT(g4273)
INPUT(g1389)
INPUT(g1706)
INPUT(g5835)
INPUT(g1171)
INPUT(g4269)
INPUT(g2399)
INPUT(g3372)
INPUT(g4983)
INPUT(g5611)
INPUT(g3618)
INPUT(g4572)
INPUT(g3143)
INPUT(g2898)
INPUT(g3343)
INPUT(g3235)
INPUT(g4543)
INPUT(g3566)
INPUT(g4534)
INPUT(g4961)
INPUT(g6398)
INPUT(g4927)
INPUT(g2259)
INPUT(g2819)
INPUT(g4414)
INPUT(g5802)
INPUT(g2852)
INPUT(g417)
INPUT(g681)
INPUT(g437)
INPUT(g351)
INPUT(g5901)
INPUT(g2886)
INPUT(g3494)
INPUT(g5511)
INPUT(g3518)
INPUT(g1604)
INPUT(g4135)
INPUT(g5092)
INPUT(g4831)
INPUT(g4382)
INPUT(g6386)
INPUT(g479)
INPUT(g3965)
INPUT(g4749)
INPUT(g2008)
INPUT(g736)
INPUT(g3933)
INPUT(g222)
INPUT(g3050)
INPUT(g5736)
INPUT(g1052)
INPUT(g58)
INPUT(g5623)
INPUT(g2122)
INPUT(g2465)
INPUT(g6483)
INPUT(g5889)
INPUT(g4495)
INPUT(g365)
INPUT(g4653)
INPUT(g3179)
INPUT(g1728)
INPUT(g2433)
INPUT(g3835)
INPUT(g6187)
INPUT(g4917)
INPUT(g1070)
INPUT(g822)
INPUT(g6027)
INPUT(g914)
INPUT(g5339)
INPUT(g4164)
INPUT(g969)
INPUT(g2807)
INPUT(g5424)
INPUT(g4054)
INPUT(g6191)
INPUT(g5077)
INPUT(g5523)
INPUT(g3680)
INPUT(g6637)
INPUT(g174)
INPUT(g1682)
INPUT(g355)
INPUT(g1087)
INPUT(g1105)
INPUT(g2342)
INPUT(g6307)
INPUT(g3802)
INPUT(g6159)
INPUT(g2255)
INPUT(g2815)
INPUT(g911)
INPUT(g43)
INPUT(g4012)
INPUT(g1748)
INPUT(g5551)
INPUT(g5742)
INPUT(g3558)
INPUT(g5499)
INPUT(g2960)
INPUT(g3901)
INPUT(g4888)
INPUT(g6251)
INPUT(g6315)
INPUT(g1373)
INPUT(g3092)
INPUT(g157)
INPUT(g2783)
INPUT(g4281)
INPUT(g3574)
INPUT(g2112)
INPUT(g1283)
INPUT(g433)
INPUT(g4297)
INPUT(g5983)
INPUT(g1459)
INPUT(g758)
INPUT(g5712)
INPUT(g4138)
INPUT(g4639)
INPUT(g6537)
INPUT(g5543)
INPUT(g1582)
INPUT(g3736)
INPUT(g5961)
INPUT(g6243)
INPUT(g632)
INPUT(g1227)
INPUT(g3889)
INPUT(g3476)
INPUT(g1664)
INPUT(g1246)
INPUT(g6128)
INPUT(g6629)
INPUT(g246)
INPUT(g4049)
INPUT(g4449)
INPUT(g2932)
INPUT(g4575)
INPUT(g4098)
INPUT(g4498)
INPUT(g528)
INPUT(g5436)
INPUT(g16)
INPUT(g3139)
INPUT(g102)
INPUT(g4584)
INPUT(g142)
INPUT(g5335)
INPUT(g5831)
INPUT(g239)
INPUT(g1216)
INPUT(g2848)
INPUT(g5805)
INPUT(g5022)
INPUT(g4019)
INPUT(g1030)
INPUT(g3672)
INPUT(g3231)
INPUT(g6490)
INPUT(g1430)
INPUT(g4452)
INPUT(g2241)
INPUT(g1564)
INPUT(g5798)
INPUT(g6148)
INPUT(g6649)
INPUT(g110)
INPUT(g884)
INPUT(g3742)
INPUT(g225)
INPUT(g4486)
INPUT(g4504)
INPUT(g5873)
INPUT(g5037)
INPUT(g2319)
INPUT(g5495)
INPUT(g4185)
INPUT(g5208)
INPUT(g2152)
INPUT(g5579)
INPUT(g5869)
INPUT(g5719)
INPUT(g1589)
INPUT(g5752)
INPUT(g6279)
INPUT(g5917)
INPUT(g2975)
INPUT(g6167)
INPUT(g3983)
INPUT(g2599)
INPUT(g1448)
INPUT(g881)
INPUT(g3712)
INPUT(g2370)
INPUT(g5164)
INPUT(g1333)
INPUT(g153)
INPUT(g6549)
INPUT(g4087)
INPUT(g4801)
INPUT(g2984)
INPUT(g3961)
INPUT(g5770)
INPUT(g962)
INPUT(g101)
INPUT(g4226)
INPUT(g6625)
INPUT(g51)
INPUT(g1018)
INPUT(g1418)
INPUT(g4045)
INPUT(g1467)
INPUT(g2461)
INPUT(g5706)
INPUT(g457)
INPUT(g2756)
INPUT(g5990)
INPUT(g471)
INPUT(g1256)
INPUT(g5029)
INPUT(g6519)
INPUT(g4169)
INPUT(g1816)
INPUT(g4369)
INPUT(g3436)
INPUT(g5787)
INPUT(g4578)
INPUT(g4459)
INPUT(g3831)
INPUT(g2514)
INPUT(g3288)
INPUT(g2403)
INPUT(g2145)
INPUT(g1700)
INPUT(g513)
INPUT(g2841)
INPUT(g5297)
INPUT(g3805)
INPUT(g2763)
INPUT(g4793)
INPUT(g952)
INPUT(g1263)
INPUT(g1950)
INPUT(g5138)
INPUT(g2307)
INPUT(g5109)
INPUT(g5791)
INPUT(g3798)
INPUT(g4664)
INPUT(g2223)
INPUT(g5808)
INPUT(g6645)
INPUT(g2016)
INPUT(g5759)
INPUT(g3873)
INPUT(g3632)
INPUT(g2315)
INPUT(g2811)
INPUT(g5957)
INPUT(g2047)
INPUT(g3869)
INPUT(g6358)
INPUT(g3719)
INPUT(g5575)
INPUT(g46)
INPUT(g3752)
INPUT(g3917)
INPUT(g4188)
INPUT(g1585)
INPUT(g4388)
INPUT(g6275)
INPUT(g6311)
INPUT(g4216)
INPUT(g1041)
INPUT(g2595)
INPUT(g2537)
INPUT(g136)
INPUT(g4430)
INPUT(g4564)
INPUT(g3454)
INPUT(g4826)
INPUT(g6239)
INPUT(g3770)
INPUT(g232)
INPUT(g5268)
INPUT(g6545)
INPUT(g2417)
INPUT(g1772)
INPUT(g4741)
INPUT(g5052)
INPUT(g5452)
INPUT(g1890)
INPUT(g2629)
INPUT(g572)
INPUT(g2130)
INPUT(g4108)
INPUT(g4308)
INPUT(g475)
INPUT(g990)
INPUT(g31)
INPUT(g3412)
INPUT(g45)
INPUT(g799)
INPUT(g3706)
INPUT(g3990)
INPUT(g5385)
INPUT(g5881)
INPUT(g1992)
INPUT(g3029)
INPUT(g3171)
INPUT(g3787)
INPUT(g812)
INPUT(g832)
INPUT(g5897)
INPUT(g4165)
INPUT(g4571)
INPUT(g3281)
INPUT(g4455)
INPUT(g2902)
INPUT(g333)
INPUT(g168)
INPUT(g2823)
INPUT(g3684)
INPUT(g3639)
INPUT(g5331)
INPUT(g3338)
INPUT(g5406)
INPUT(g3791)
INPUT(g269)
INPUT(g401)
INPUT(g6040)
INPUT(g441)
INPUT(g5105)
INPUT(g3808)
INPUT(g9)
INPUT(g3759)
INPUT(g4467)
INPUT(g3957)
INPUT(g4093)
INPUT(g1760)
INPUT(g6151)
INPUT(g6351)
INPUT(g160)
INPUT(g5445)
INPUT(g5373)
INPUT(g2279)
INPUT(g3498)
INPUT(g586)
INPUT(g869)
INPUT(g2619)
INPUT(g1183)
INPUT(g1608)
INPUT(g4197)
INPUT(g5283)
INPUT(g1779)
INPUT(g2652)
INPUT(g5459)
INPUT(g2193)
INPUT(g2393)
INPUT(g5767)
INPUT(g661)
INPUT(g4950)
INPUT(g5535)
INPUT(g2834)
INPUT(g1361)
INPUT(g3419)
INPUT(g6235)
INPUT(g1146)
INPUT(g2625)
INPUT(g150)
INPUT(g1696)
INPUT(g6555)
INPUT(g859)
INPUT(g3385)
INPUT(g3881)
INPUT(g6621)
INPUT(g3470)
INPUT(g3897)
INPUT(g518)
INPUT(g3025)
INPUT(g538)
INPUT(g2606)
INPUT(g1472)
INPUT(g6113)
INPUT(g542)
INPUT(g5188)
INPUT(g5689)
INPUT(g1116)
INPUT(g405)
INPUT(g5216)
INPUT(g6494)
INPUT(g4669)
INPUT(g5428)
INPUT(g996)
INPUT(g4531)
INPUT(g2860)
INPUT(g4743)
INPUT(g6593)
INPUT(g2710)
INPUT(g215)
INPUT(g4411)
INPUT(g1413)
INPUT(g4474)
INPUT(g5308)
INPUT(g6641)
INPUT(g3045)
INPUT(g6)
INPUT(g1936)
INPUT(g55)
INPUT(g504)
INPUT(g2587)
INPUT(g4480)
INPUT(g2311)
INPUT(g3602)
INPUT(g5571)
INPUT(g3578)
INPUT(g468)
INPUT(g5448)
INPUT(g3767)
INPUT(g5827)
INPUT(g3582)
INPUT(g6271)
INPUT(g4688)
INPUT(g5774)
INPUT(g2380)
INPUT(g5196)
INPUT(g5396)
INPUT(g3227)
INPUT(g2020)
INPUT(g4000)
INPUT(g1079)
INPUT(g6541)
INPUT(g3203)
INPUT(g1668)
INPUT(g4760)
INPUT(g262)
INPUT(g1840)
INPUT(g70)
INPUT(g5467)
INPUT(g460)
INPUT(g6209)
INPUT(g74)
INPUT(g5290)
INPUT(g655)
INPUT(g3502)
INPUT(g2204)
INPUT(g5256)
INPUT(g4608)
INPUT(g794)
INPUT(g4023)
INPUT(g4423)
INPUT(g3689)
INPUT(g5381)
INPUT(g5685)
INPUT(g703)
INPUT(g5421)
INPUT(g862)
INPUT(g3247)
INPUT(g2040)
INPUT(g4999)
INPUT(g4146)
INPUT(g4633)
INPUT(g1157)
INPUT(g5723)
INPUT(g4732)
INPUT(g5101)
INPUT(g5817)
INPUT(g2151)
INPUT(g2351)
INPUT(g2648)
INPUT(g6736)
INPUT(g4944)
INPUT(g4072)
INPUT(g344)
INPUT(g4443)
INPUT(g3466)
INPUT(g4116)
INPUT(g5041)
INPUT(g5441)
INPUT(g4434)
INPUT(g3827)
INPUT(g6500)
INPUT(g5673)
INPUT(g3133)
INPUT(g3333)
INPUT(g979)
INPUT(g4681)
INPUT(g298)
INPUT(g3774)
INPUT(g2667)
INPUT(g3396)
INPUT(g4210)
INPUT(g1894)
INPUT(g2988)
INPUT(g3538)
INPUT(g301)
INPUT(g341)
INPUT(g827)
INPUT(g1075)
INPUT(g6077)
INPUT(g2555)
INPUT(g5011)
INPUT(g199)
INPUT(g6523)
INPUT(g1526)
INPUT(g4601)
INPUT(g854)
INPUT(g1484)
INPUT(g4922)
INPUT(g5080)
INPUT(g5863)
INPUT(g4581)
INPUT(g3021)
INPUT(g2518)
INPUT(g2567)
INPUT(g568)
INPUT(g3263)
INPUT(g6613)
INPUT(g6044)
INPUT(g6444)
INPUT(g2965)
INPUT(g5857)
INPUT(g1616)
INPUT(g890)
INPUT(g5976)
INPUT(g3562)
INPUT(g4294)
INPUT(g1404)
INPUT(g3723)
INPUT(g3817)
INPUT(g93)
INPUT(g4501)
INPUT(g287)
INPUT(g2724)
INPUT(g4704)
INPUT(g22)
INPUT(g2878)
INPUT(g5220)
INPUT(g617)
INPUT(g637)
INPUT(g316)
INPUT(g1277)
INPUT(g6513)
INPUT(g336)
INPUT(g2882)
INPUT(g933)
INPUT(g1906)
INPUT(g305)
INPUT(g8)
INPUT(g3368)
INPUT(g2799)
INPUT(g887)
INPUT(g5327)
INPUT(g4912)
INPUT(g4157)
INPUT(g2541)
INPUT(g2153)
INPUT(g550)
INPUT(g255)
INPUT(g1945)
INPUT(g5240)
INPUT(g1478)
INPUT(g3080)
INPUT(g3863)
INPUT(g1959)
INPUT(g3480)
INPUT(g6653)
INPUT(g6719)
INPUT(g2864)
INPUT(g4894)
INPUT(g5681)
INPUT(g3857)
INPUT(g3976)
INPUT(g499)
INPUT(g5413)
INPUT(g1002)
INPUT(g776)
INPUT(g28)
INPUT(g1236)
INPUT(g4646)
INPUT(g2476)
INPUT(g1657)
INPUT(g2375)
INPUT(g63)
INPUT(g6012)
INPUT(g358)
INPUT(g896)
INPUT(g967)
INPUT(g3423)
INPUT(g283)
INPUT(g3161)
INPUT(g2384)
INPUT(g3361)
INPUT(g6675)
INPUT(g4616)
INPUT(g4561)
INPUT(g2024)
INPUT(g3451)
INPUT(g2795)
INPUT(g613)
INPUT(g4527)
INPUT(g1844)
INPUT(g5937)
INPUT(g4546)
INPUT(g3103)
INPUT(g2523)
INPUT(g3303)
INPUT(g2643)
INPUT(g6109)
INPUT(g1489)
INPUT(g5390)
INPUT(g194)
INPUT(g2551)
INPUT(g5156)
INPUT(g3072)
INPUT(g1242)
INPUT(g47)
INPUT(g3443)
INPUT(g4277)
INPUT(g1955)
INPUT(g6049)
INPUT(g3034)
INPUT(g2273)
INPUT(g6715)
INPUT(g4771)
INPUT(g6098)
INPUT(g3147)
INPUT(g3347)
INPUT(g2269)
INPUT(g191)
INPUT(g2712)
INPUT(g626)
INPUT(g2729)
INPUT(g5357)
INPUT(g4991)
INPUT(g6019)
INPUT(g4709)
INPUT(g6419)
INPUT(g6052)
INPUT(g2927)
INPUT(g4340)
INPUT(g5929)
INPUT(g4907)
INPUT(g3317)
INPUT(g4035)
INPUT(g2946)
INPUT(g918)
INPUT(g4082)
INPUT(g6486)
INPUT(g2036)
INPUT(g577)
INPUT(g1620)
INPUT(g2831)
INPUT(g667)
INPUT(g930)
INPUT(g3937)
INPUT(g5782)
INPUT(g817)
INPUT(g1249)
INPUT(g837)
INPUT(g3668)
INPUT(g599)
INPUT(g5475)
INPUT(g739)
INPUT(g5949)
INPUT(g6682)
INPUT(g6105)
INPUT(g904)
INPUT(g2873)
INPUT(g1854)
INPUT(g5084)
INPUT(g5603)
INPUT(g4222)
INPUT(g2495)
INPUT(g2437)
INPUT(g2102)
INPUT(g2208)
INPUT(g2579)
INPUT(g4064)
INPUT(g4899)
INPUT(g2719)
INPUT(g4785)
INPUT(g5583)
INPUT(g781)
INPUT(g6173)
INPUT(g6373)
INPUT(g2917)
INPUT(g686)
INPUT(g1252)
INPUT(g671)
INPUT(g2265)
INPUT(g6283)
INPUT(g6369)
INPUT(g5276)
INPUT(g6459)
INPUT(g901)
INPUT(g4194)
INPUT(g5527)
INPUT(g4489)
INPUT(g1974)
INPUT(g1270)
INPUT(g4966)
INPUT(g6415)
INPUT(g6227)
INPUT(g3929)
INPUT(g5503)
INPUT(g4242)
INPUT(g5925)
INPUT(g1124)
INPUT(g4955)
INPUT(g5224)
INPUT(g2012)
INPUT(g6203)
INPUT(g5120)
INPUT(g5320)
INPUT(g2389)
INPUT(g4438)
INPUT(g2429)
INPUT(g2787)
INPUT(g1287)
INPUT(g2675)
INPUT(g66)
INPUT(g4836)
INPUT(g1199)
INPUT(g1399)
INPUT(g5547)
INPUT(g3782)
INPUT(g6428)
INPUT(g2138)
INPUT(g3661)
INPUT(g2338)
INPUT(g4229)
INPUT(g6247)
INPUT(g2791)
INPUT(g3949)
INPUT(g1291)
INPUT(g5945)
INPUT(g5244)
INPUT(g2759)
INPUT(g6741)
INPUT(g785)
INPUT(g1259)
INPUT(g3484)
INPUT(g209)
INPUT(g6609)
INPUT(g5517)
INPUT(g2449)
INPUT(g2575)
INPUT(g65)
INPUT(g2715)
INPUT(g936)
INPUT(g2098)
INPUT(g4462)
INPUT(g604)
INPUT(g6589)
INPUT(g1886)
INPUT(g6466)
INPUT(g6365)
INPUT(g6711)
INPUT(g429)
INPUT(g1870)
INPUT(g4249)
INPUT(g6455)
INPUT(g3004)
INPUT(g1825)
INPUT(g6133)
INPUT(g1008)
INPUT(g4392)
INPUT(g5002)
INPUT(g3546)
INPUT(g5236)
INPUT(g1768)
INPUT(g4854)
INPUT(g3925)
INPUT(g6509)
INPUT(g732)
INPUT(g2504)
INPUT(g1322)
INPUT(g4520)
INPUT(g4219)
INPUT(g2185)
INPUT(g37)
INPUT(g4031)
INPUT(g2070)
INPUT(g4812)
INPUT(g6093)
INPUT(g968)
INPUT(g4176)
INPUT(g4005)
INPUT(g4405)
INPUT(g872)
INPUT(g6181)
INPUT(g6381)
INPUT(g4765)
INPUT(g5563)
INPUT(g1395)
INPUT(g1913)
INPUT(g2331)
INPUT(g6263)
INPUT(g50)
INPUT(g3945)
INPUT(g347)
INPUT(g5731)
INPUT(g4473)
INPUT(g1266)
INPUT(g5489)
INPUT(g714)
INPUT(g2748)
INPUT(g5471)
INPUT(g4540)
INPUT(g6723)
INPUT(g6605)
INPUT(g2445)
INPUT(g2173)
INPUT(g4287)
INPUT(g2491)
INPUT(g4849)
INPUT(g2169)
INPUT(g2283)
INPUT(g6585)
INPUT(g121)
INPUT(g2407)
INPUT(g2868)
INPUT(g2767)
INPUT(g1783)
INPUT(g3310)
INPUT(g1312)
INPUT(g5212)
INPUT(g4245)
INPUT(g645)
INPUT(g4291)
INPUT(g79)
INPUT(g182)
INPUT(g1129)
INPUT(g2227)
INPUT(g6058)
INPUT(g4207)
INPUT(g2246)
INPUT(g1830)
INPUT(g3590)
INPUT(g392)
INPUT(g1592)
INPUT(g6505)
INPUT(g6411)
INPUT(g1221)
INPUT(g5921)
INPUT(g106)
INPUT(g146)
INPUT(g218)
INPUT(g6474)
INPUT(g1932)
INPUT(g1624)
INPUT(g5062)
INPUT(g5462)
INPUT(g2689)
INPUT(g6573)
INPUT(g1677)
INPUT(g2028)
INPUT(g2671)
INPUT(g1576)
INPUT(g4408)
INPUT(g34)
INPUT(g1848)
INPUT(g3089)
INPUT(g3731)
INPUT(g86)
INPUT(g5485)
INPUT(g2741)
INPUT(g802)
INPUT(g2638)
INPUT(g4122)
INPUT(g4322)
INPUT(g5941)
INPUT(g2108)
INPUT(g6000)
INPUT(g25)
INPUT(g1644)
INPUT(g595)
INPUT(g2217)
INPUT(g1319)
INPUT(g2066)
INPUT(g1152)
INPUT(g5252)
INPUT(g2165)
INPUT(g2571)
INPUT(g5176)
INPUT(g391)
INPUT(g5005)
INPUT(g2711)
INPUT(g6023)
INPUT(g1211)
INPUT(g2827)
INPUT(g6423)
INPUT(g875)
INPUT(g4859)
INPUT(g424)
INPUT(g1274)
INPUT(g1426)
INPUT(g85)
INPUT(g2803)
INPUT(g6451)
INPUT(g1821)
INPUT(g2509)
INPUT(g5073)
INPUT(g1280)
INPUT(g4815)
INPUT(g6346)
INPUT(g6633)
INPUT(g5124)
INPUT(g1083)
INPUT(g6303)
INPUT(g5069)
INPUT(g2994)
INPUT(g650)
INPUT(g1636)
INPUT(g3921)
INPUT(g2093)
INPUT(g6732)
INPUT(g1306)
INPUT(g5377)
INPUT(g1061)
INPUT(g3462)
INPUT(g2181)
INPUT(g956)
INPUT(g1756)
INPUT(g5849)
INPUT(g4112)
INPUT(g2685)
INPUT(g2197)
INPUT(g6116)
INPUT(g2421)
INPUT(g1046)
INPUT(g482)
INPUT(g4401)
INPUT(g6434)
INPUT(g1514)
INPUT(g329)
INPUT(g6565)
INPUT(g2950)
INPUT(g4129)
INPUT(g1345)
INPUT(g6533)
INPUT(g3298)
INPUT(g3085)
INPUT(g4727)
INPUT(g6697)
INPUT(g1536)
INPUT(g3941)
INPUT(g370)
INPUT(g5694)
INPUT(g1858)
INPUT(g446)
INPUT(g4932)
INPUT(g3219)
INPUT(g1811)
INPUT(g3431)
INPUT(g6601)
INPUT(g3376)
INPUT(g2441)
INPUT(g1874)
INPUT(g4349)
INPUT(g6581)
INPUT(g6597)
INPUT(g5008)
INPUT(g3610)
INPUT(g2890)
INPUT(g1978)
INPUT(g1612)
INPUT(g112)
INPUT(g2856)
INPUT(g6479)
INPUT(g1982)
INPUT(g6668)
INPUT(g5228)
INPUT(g4119)
INPUT(g6390)
INPUT(g1542)
INPUT(g4258)
INPUT(g4818)
INPUT(g5033)
INPUT(g4717)
INPUT(g1554)
INPUT(g3849)
INPUT(g6704)
INPUT(g3199)
INPUT(g5845)
INPUT(g4975)
INPUT(g790)
INPUT(g5913)
INPUT(g1902)
INPUT(g6163)
INPUT(g4125)
INPUT(g4821)
INPUT(g4939)
INPUT(g1056)
INPUT(g3207)
INPUT(g4483)
INPUT(g3259)
INPUT(g5142)
INPUT(g5248)
INPUT(g2126)
INPUT(g3694)
INPUT(g5481)
INPUT(g1964)
INPUT(g5097)
INPUT(g3215)
INPUT(g4027)
INPUT(g111)
INPUT(g4427)
INPUT(g7)
INPUT(g2779)
INPUT(g4200)
INPUT(g4446)
INPUT(g1720)
INPUT(g1367)
INPUT(g5112)
INPUT(g19)
INPUT(g4145)
INPUT(g2161)
INPUT(g376)
INPUT(g2361)
INPUT(g4191)
INPUT(g582)
INPUT(g2051)
INPUT(g1193)
INPUT(g5401)
INPUT(g3408)
INPUT(g2327)
INPUT(g907)
INPUT(g947)
INPUT(g1834)
INPUT(g3594)
INPUT(g2999)
INPUT(g5727)
INPUT(g2303)
INPUT(g6661)
INPUT(g3065)
INPUT(g699)
INPUT(g723)
INPUT(g5703)
INPUT(g546)
INPUT(g2472)
INPUT(g5953)
INPUT(g3096)
INPUT(g6439)
INPUT(g1740)
INPUT(g3550)
INPUT(g3845)
INPUT(g2116)
INPUT(g5677)
INPUT(g3195)
INPUT(g3913)
INPUT(g4537)
INPUT(g1687)
INPUT(g2681)
INPUT(g2533)
INPUT(g324)
INPUT(g2697)
INPUT(g5747)
INPUT(g4417)
INPUT(g6561)
INPUT(g1141)
INPUT(g1570)
INPUT(g2413)
INPUT(g1710)
INPUT(g6527)
INPUT(g6404)
INPUT(g3255)
INPUT(g1691)
INPUT(g2936)
INPUT(g5644)
INPUT(g5152)
INPUT(g5352)
INPUT(g4213)
INPUT(g6120)
INPUT(g2775)
INPUT(g2922)
INPUT(g1111)
INPUT(g5893)
INPUT(g1311)
INPUT(g3267)
INPUT(g6617)
INPUT(g2060)
INPUT(g4512)
INPUT(g5599)
INPUT(g3401)
INPUT(g4366)
INPUT(g3676)
INPUT(g94)
INPUT(g3129)
INPUT(g3329)
INPUT(g5170)
INPUT(g4456)
INPUT(g5821)
INPUT(g6299)
INPUT(g1239)
INPUT(g3727)
INPUT(g2079)
INPUT(g4698)
INPUT(g3703)
INPUT(g1559)
INPUT(g943)
INPUT(g411)
INPUT(g6140)
INPUT(g3953)
INPUT(g3068)
INPUT(g2704)
INPUT(g6035)
INPUT(g6082)
INPUT(g49)
INPUT(g1300)
INPUT(g4057)
INPUT(g5200)
INPUT(g4843)
INPUT(g5046)
INPUT(g2250)
INPUT(g319)
INPUT(g4549)
INPUT(g2453)
INPUT(g5841)
INPUT(g5763)
INPUT(g3747)
INPUT(g5637)
INPUT(g2912)
INPUT(g2357)
INPUT(g4232)
INPUT(g164)
INPUT(g4253)
INPUT(g5016)
INPUT(g3119)
INPUT(g1351)
INPUT(g1648)
INPUT(g4519)
INPUT(g5115)
INPUT(g3352)
INPUT(g6657)
INPUT(g4552)
INPUT(g3893)
INPUT(g3211)
INPUT(g5654)
INPUT(g929)
INPUT(g3274)
INPUT(g5595)
INPUT(g3614)
INPUT(g2894)
INPUT(g3125)
INPUT(g3325)
INPUT(g3821)
INPUT(g4141)
INPUT(g4570)
INPUT(g5272)
INPUT(g2735)
INPUT(g728)
INPUT(g6295)
INPUT(g5417)
INPUT(g2661)
INPUT(g1988)
INPUT(g5128)
INPUT(g1548)
INPUT(g3106)
INPUT(g4659)
INPUT(g4358)
INPUT(g1792)
INPUT(g2084)
INPUT(g3061)
INPUT(g3187)
INPUT(g4311)
INPUT(g2583)
INPUT(g3003)
INPUT(g1094)
INPUT(g3841)
INPUT(g4284)
INPUT(g3763)
INPUT(g3191)
INPUT(g4239)
INPUT(g3391)
INPUT(g4180)
INPUT(g691)
INPUT(g534)
INPUT(g5366)
INPUT(g385)
INPUT(g2004)
INPUT(g2527)
INPUT(g5456)
INPUT(g4420)
INPUT(g5148)
INPUT(g4507)
INPUT(g5348)
INPUT(g3223)
INPUT(g4931)
INPUT(g2970)
INPUT(g5698)
INPUT(g3416)
INPUT(g5260)
INPUT(g1521)
INPUT(g3522)
INPUT(g3115)
INPUT(g3251)
INPUT(g1)
INPUT(g4628)
INPUT(g1996)
INPUT(g3447)
INPUT(g4515)
INPUT(g4204)
INPUT(g4300)
INPUT(g1724)
INPUT(g1379)
INPUT(g3654)
INPUT(g12)
INPUT(g1878)
INPUT(g5619)
INPUT(g71)
INPUT(g59)
OUTPUT(g7243)
OUTPUT(g7245)
OUTPUT(g7257)
OUTPUT(g7260)
OUTPUT(g7540)
OUTPUT(g7916)
OUTPUT(g7946)
OUTPUT(g8132)
OUTPUT(g8178)
OUTPUT(g8215)
OUTPUT(g8235)
OUTPUT(g8277)
OUTPUT(g8279)
OUTPUT(g8283)
OUTPUT(g8291)
OUTPUT(g8342)
OUTPUT(g8344)
OUTPUT(g8353)
OUTPUT(g8358)
OUTPUT(g8398)
OUTPUT(g8403)
OUTPUT(g8416)
OUTPUT(g8475)
OUTPUT(g8719)
OUTPUT(g8783)
OUTPUT(g8784)
OUTPUT(g8785)
OUTPUT(g8786)
OUTPUT(g8787)
OUTPUT(g8788)
OUTPUT(g8789)
OUTPUT(g8839)
OUTPUT(g8870)
OUTPUT(g8915)
OUTPUT(g8916)
OUTPUT(g8917)
OUTPUT(g8918)
OUTPUT(g8919)
OUTPUT(g8920)
OUTPUT(g9019)
OUTPUT(g9048)
OUTPUT(g9251)
OUTPUT(g9497)
OUTPUT(g9553)
OUTPUT(g9555)
OUTPUT(g9615)
OUTPUT(g9617)
OUTPUT(g9680)
OUTPUT(g9682)
OUTPUT(g9741)
OUTPUT(g9743)
OUTPUT(g9817)
OUTPUT(g10122)
OUTPUT(g10306)
OUTPUT(g10500)
OUTPUT(g10527)
OUTPUT(g11349)
OUTPUT(g11388)
OUTPUT(g11418)
OUTPUT(g11447)
OUTPUT(g11678)
OUTPUT(g11770)
OUTPUT(g12184)
OUTPUT(g12238)
OUTPUT(g12300)
OUTPUT(g12350)
OUTPUT(g12368)
OUTPUT(g12422)
OUTPUT(g12470)
OUTPUT(g12832)
OUTPUT(g12919)
OUTPUT(g12923)
OUTPUT(g13039)
OUTPUT(g13049)
OUTPUT(g13068)
OUTPUT(g13085)
OUTPUT(g13099)
OUTPUT(g13259)
OUTPUT(g13272)
OUTPUT(g13865)
OUTPUT(g13881)
OUTPUT(g13895)
OUTPUT(g13906)
OUTPUT(g13926)
OUTPUT(g13966)
OUTPUT(g14096)
OUTPUT(g14125)
OUTPUT(g14147)
OUTPUT(g14167)
OUTPUT(g14189)
OUTPUT(g14201)
OUTPUT(g14217)
OUTPUT(g14421)
OUTPUT(g14451)
OUTPUT(g14518)
OUTPUT(g14597)
OUTPUT(g14635)
OUTPUT(g14662)
OUTPUT(g14673)
OUTPUT(g14694)
OUTPUT(g14705)
OUTPUT(g14738)
OUTPUT(g14749)
OUTPUT(g14779)
OUTPUT(g14828)
OUTPUT(g16603)
OUTPUT(g16624)
OUTPUT(g16627)
OUTPUT(g16656)
OUTPUT(g16659)
OUTPUT(g16686)
OUTPUT(g16693)
OUTPUT(g16718)
OUTPUT(g16722)
OUTPUT(g16744)
OUTPUT(g16748)
OUTPUT(g16775)
OUTPUT(g16874)
OUTPUT(g16924)
OUTPUT(g16955)
OUTPUT(g17291)
OUTPUT(g17316)
OUTPUT(g17320)
OUTPUT(g17400)
OUTPUT(g17404)
OUTPUT(g17423)
OUTPUT(g17519)
OUTPUT(g17577)
OUTPUT(g17580)
OUTPUT(g17604)
OUTPUT(g17607)
OUTPUT(g17639)
OUTPUT(g17646)
OUTPUT(g17649)
OUTPUT(g17674)
OUTPUT(g17678)
OUTPUT(g17685)
OUTPUT(g17688)
OUTPUT(g17711)
OUTPUT(g17715)
OUTPUT(g17722)
OUTPUT(g17739)
OUTPUT(g17743)
OUTPUT(g17760)
OUTPUT(g17764)
OUTPUT(g17778)
OUTPUT(g17787)
OUTPUT(g17813)
OUTPUT(g17819)
OUTPUT(g17845)
OUTPUT(g17871)
OUTPUT(g18092)
OUTPUT(g18094)
OUTPUT(g18095)
OUTPUT(g18096)
OUTPUT(g18097)
OUTPUT(g18098)
OUTPUT(g18099)
OUTPUT(g18100)
OUTPUT(g18101)
OUTPUT(g18881)
OUTPUT(g19334)
OUTPUT(g19357)
OUTPUT(g20049)
OUTPUT(g20557)
OUTPUT(g20652)
OUTPUT(g20654)
OUTPUT(g20763)
OUTPUT(g20899)
OUTPUT(g20901)
OUTPUT(g21176)
OUTPUT(g21245)
OUTPUT(g21270)
OUTPUT(g21292)
OUTPUT(g21698)
OUTPUT(g21727)
OUTPUT(g23002)
OUTPUT(g23190)
OUTPUT(g23612)
OUTPUT(g23652)
OUTPUT(g23683)
OUTPUT(g23759)
OUTPUT(g24151)
OUTPUT(g25114)
OUTPUT(g25167)
OUTPUT(g25219)
OUTPUT(g25259)
OUTPUT(g25582)
OUTPUT(g25583)
OUTPUT(g25584)
OUTPUT(g25585)
OUTPUT(g25586)
OUTPUT(g25587)
OUTPUT(g25588)
OUTPUT(g25589)
OUTPUT(g25590)
OUTPUT(g26801)
OUTPUT(g26875)
OUTPUT(g26876)
OUTPUT(g26877)
OUTPUT(g27831)
OUTPUT(g28030)
OUTPUT(g28041)
OUTPUT(g28042)
OUTPUT(g28753)
OUTPUT(g29210)
OUTPUT(g29211)
OUTPUT(g29212)
OUTPUT(g29213)
OUTPUT(g29214)
OUTPUT(g29215)
OUTPUT(g29216)
OUTPUT(g29217)
OUTPUT(g29218)
OUTPUT(g29219)
OUTPUT(g29220)
OUTPUT(g29221)
OUTPUT(g30327)
OUTPUT(g30329)
OUTPUT(g30330)
OUTPUT(g30331)
OUTPUT(g30332)
OUTPUT(g31521)
OUTPUT(g31656)
OUTPUT(g31665)
OUTPUT(g31793)
OUTPUT(g31860)
OUTPUT(g31861)
OUTPUT(g31862)
OUTPUT(g31863)
OUTPUT(g32185)
OUTPUT(g32429)
OUTPUT(g32454)
OUTPUT(g32975)
OUTPUT(g33079)
OUTPUT(g33435)
OUTPUT(g33533)
OUTPUT(g33636)
OUTPUT(g33659)
OUTPUT(g33874)
OUTPUT(g33894)
OUTPUT(g33935)
OUTPUT(g33945)
OUTPUT(g33946)
OUTPUT(g33947)
OUTPUT(g33948)
OUTPUT(g33949)
OUTPUT(g33950)
OUTPUT(g33959)
OUTPUT(g34201)
OUTPUT(g34221)
OUTPUT(g34232)
OUTPUT(g34233)
OUTPUT(g34234)
OUTPUT(g34235)
OUTPUT(g34236)
OUTPUT(g34237)
OUTPUT(g34238)
OUTPUT(g34239)
OUTPUT(g34240)
OUTPUT(g34383)
OUTPUT(g34425)
OUTPUT(g34435)
OUTPUT(g34436)
OUTPUT(g34437)
OUTPUT(g34597)
OUTPUT(g34788)
OUTPUT(g34839)
OUTPUT(g34913)
OUTPUT(g34915)
OUTPUT(g34917)
OUTPUT(g34919)
OUTPUT(g34921)
OUTPUT(g34923)
OUTPUT(g34925)
OUTPUT(g34927)
OUTPUT(g34956)
OUTPUT(g34972)
OUTPUT(g24168)
OUTPUT(g24178)
OUTPUT(g12833)
OUTPUT(g24174)
OUTPUT(g24181)
OUTPUT(g24172)
OUTPUT(g24161)
OUTPUT(g24177)
OUTPUT(g24171)
OUTPUT(g24163)
OUTPUT(g24170)
OUTPUT(g24185)
OUTPUT(g24164)
OUTPUT(g24173)
OUTPUT(g24162)
OUTPUT(g24179)
OUTPUT(g24180)
OUTPUT(g24175)
OUTPUT(g24183)
OUTPUT(g24166)
OUTPUT(g24176)
OUTPUT(g24184)
OUTPUT(g24169)
OUTPUT(g24182)
OUTPUT(g24165)
OUTPUT(g24167)
OUTPUT(g33046)
OUTPUT(g34441)
OUTPUT(g33982)
OUTPUT(g25751)
OUTPUT(g34007)
OUTPUT(g24276)
OUTPUT(g30381)
OUTPUT(g640)
OUTPUT(g31877)
OUTPUT(g30405)
OUTPUT(g25604)
OUTPUT(g25607)
OUTPUT(g30416)
OUTPUT(g30466)
OUTPUT(g25736)
OUTPUT(g34617)
OUTPUT(g33974)
OUTPUT(g30505)
OUTPUT(g33554)
OUTPUT(g30432)
OUTPUT(g33064)
OUTPUT(g34881)
OUTPUT(g6027)
OUTPUT(g24216)
OUTPUT(g24232)
OUTPUT(g34733)
OUTPUT(g34882)
OUTPUT(g33026)
OUTPUT(g31867)
OUTPUT(g25668)
OUTPUT(g24344)
OUTPUT(g4232)
OUTPUT(g33966)
OUTPUT(g33550)
OUTPUT(g3625)
OUTPUT(g30393)
OUTPUT(g31880)
OUTPUT(g29248)
OUTPUT(g4571)
OUTPUT(g24274)
OUTPUT(g31920)
OUTPUT(g33973)
OUTPUT(g30360)
OUTPUT(g34460)
OUTPUT(g30494)
OUTPUT(g30384)
OUTPUT(g24340)
OUTPUT(g29223)
OUTPUT(g26881)
OUTPUT(g31925)
OUTPUT(g34252)
OUTPUT(g30489)
OUTPUT(g29301)
OUTPUT(g6373)
OUTPUT(g33022)
OUTPUT(g30496)
OUTPUT(g33043)
OUTPUT(g28062)
OUTPUT(g29263)
OUTPUT(g30533)
OUTPUT(g24256)
OUTPUT(g34015)
OUTPUT(g34031)
OUTPUT(g34452)
OUTPUT(g34646)
OUTPUT(g34001)
OUTPUT(g25633)
OUTPUT(g24259)
OUTPUT(g33049)
OUTPUT(g34609)
OUTPUT(g31869)
OUTPUT(g30490)
OUTPUT(g30427)
OUTPUT(g21894)
OUTPUT(g33965)
OUTPUT(g34645)
OUTPUT(g3317)
OUTPUT(g33571)
OUTPUT(g34267)
OUTPUT(g26971)
OUTPUT(g34644)
OUTPUT(g3618)
OUTPUT(g30534)
OUTPUT(g33535)
OUTPUT(g30498)
OUTPUT(g25728)
OUTPUT(g25743)
OUTPUT(g25684)
OUTPUT(g25613)
OUTPUT(g34438)
OUTPUT(g24244)
OUTPUT(g30439)
OUTPUT(g30541)
OUTPUT(g30519)
OUTPUT(g25621)
OUTPUT(g34807)
OUTPUT(g25599)
OUTPUT(g31924)
OUTPUT(g24235)
OUTPUT(g34036)
OUTPUT(g30476)
OUTPUT(g5623)
OUTPUT(g30429)
OUTPUT(g32997)
OUTPUT(g33063)
OUTPUT(g30424)
OUTPUT(g32977)
OUTPUT(g34026)
OUTPUT(g30420)
OUTPUT(g637)
OUTPUT(g6012)
OUTPUT(g33560)
OUTPUT(g29226)
OUTPUT(g25619)
OUTPUT(g28076)
OUTPUT(g34455)
OUTPUT(g30457)
OUTPUT(g5637)
OUTPUT(g33625)
OUTPUT(g34790)
OUTPUT(g30414)
OUTPUT(g26966)
OUTPUT(g31923)
OUTPUT(g6315)
OUTPUT(g25656)
OUTPUT(g30390)
OUTPUT(g26935)
OUTPUT(g34727)
OUTPUT(g25594)
OUTPUT(g26963)
OUTPUT(g34034)
OUTPUT(g33541)
OUTPUT(g28093)
OUTPUT(g24236)
OUTPUT(g30404)
OUTPUT(g28051)
OUTPUT(g29303)
OUTPUT(g26917)
OUTPUT(g25741)
OUTPUT(g33624)
OUTPUT(g31882)
OUTPUT(g24337)
OUTPUT(g34911)
OUTPUT(g33963)
OUTPUT(g34627)
OUTPUT(g29282)
OUTPUT(g1418)
OUTPUT(g25676)
OUTPUT(g33013)
OUTPUT(g32981)
OUTPUT(g34993)
OUTPUT(g30483)
OUTPUT(g875)
OUTPUT(g32994)
OUTPUT(g28070)
OUTPUT(g34806)
OUTPUT(g30453)
OUTPUT(g33539)
OUTPUT(g30526)
OUTPUT(g26951)
OUTPUT(g34035)
OUTPUT(g34636)
OUTPUT(g32978)
OUTPUT(g6668)
OUTPUT(g30348)
OUTPUT(g24336)
OUTPUT(g3092)
OUTPUT(g24250)
OUTPUT(g6490)
OUTPUT(g29236)
OUTPUT(g29298)
OUTPUT(g1576)
OUTPUT(g30499)
OUTPUT(g33976)
OUTPUT(g32996)
OUTPUT(g30335)
OUTPUT(g31878)
OUTPUT(g34637)
OUTPUT(g25693)
OUTPUT(g30528)
OUTPUT(g25661)
OUTPUT(g4012)
OUTPUT(g24251)
OUTPUT(g30521)
OUTPUT(g26960)
OUTPUT(g24239)
OUTPUT(g34259)
OUTPUT(g30474)
OUTPUT(g6351)
OUTPUT(g33016)
OUTPUT(g34643)
OUTPUT(g31905)
OUTPUT(g30510)
OUTPUT(g29239)
OUTPUT(g26897)
OUTPUT(g34729)
OUTPUT(g34625)
OUTPUT(g34800)
OUTPUT(g24353)
OUTPUT(g33029)
OUTPUT(g21903)
OUTPUT(g33615)
OUTPUT(g24253)
OUTPUT(g24281)
OUTPUT(g33997)
OUTPUT(g25651)
OUTPUT(g34997)
OUTPUT(g34263)
OUTPUT(g24237)
OUTPUT(g33584)
OUTPUT(g24280)
OUTPUT(g26920)
OUTPUT(g33548)
OUTPUT(g29296)
OUTPUT(g30338)
OUTPUT(g21895)
OUTPUT(g33588)
OUTPUT(g31886)
OUTPUT(g34041)
OUTPUT(g30495)
OUTPUT(g3661)
OUTPUT(g29279)
OUTPUT(g25655)
OUTPUT(g34795)
OUTPUT(g24269)
OUTPUT(g30403)
OUTPUT(g33042)
OUTPUT(g30419)
OUTPUT(g34023)
OUTPUT(g28090)
OUTPUT(g31926)
OUTPUT(g34642)
OUTPUT(g30370)
OUTPUT(g34448)
OUTPUT(g26946)
OUTPUT(g5794)
OUTPUT(g34610)
OUTPUT(g24209)
OUTPUT(g28047)
OUTPUT(g24206)
OUTPUT(g26891)
OUTPUT(g30504)
OUTPUT(g34798)
OUTPUT(g25669)
OUTPUT(g30480)
OUTPUT(g33027)
OUTPUT(g33972)
OUTPUT(g28077)
OUTPUT(g25697)
OUTPUT(g28099)
OUTPUT(g26947)
OUTPUT(g24350)
OUTPUT(g24210)
OUTPUT(g30455)
OUTPUT(g28084)
OUTPUT(g33993)
OUTPUT(g802)
OUTPUT(g30444)
OUTPUT(g33537)
OUTPUT(g25650)
OUTPUT(g31915)
OUTPUT(g25625)
OUTPUT(g30328)
OUTPUT(g5666)
OUTPUT(g30366)
OUTPUT(g33593)
OUTPUT(g25755)
OUTPUT(g30502)
OUTPUT(g33036)
OUTPUT(g25595)
OUTPUT(g34462)
OUTPUT(g33024)
OUTPUT(g33552)
OUTPUT(g34014)
OUTPUT(g29273)
OUTPUT(g25748)
OUTPUT(g34638)
OUTPUT(g30341)
OUTPUT(g26899)
OUTPUT(g6023)
OUTPUT(g30336)
OUTPUT(g5335)
OUTPUT(g26940)
OUTPUT(g25622)
OUTPUT(g34447)
OUTPUT(g25709)
OUTPUT(g33613)
OUTPUT(g25749)
OUTPUT(g25704)
OUTPUT(g33053)
OUTPUT(g3676)
OUTPUT(g30555)
OUTPUT(g25601)
OUTPUT(g33971)
OUTPUT(g26892)
OUTPUT(g1083)
OUTPUT(g26915)
OUTPUT(g33008)
OUTPUT(g30538)
OUTPUT(g3794)
OUTPUT(g25750)
OUTPUT(g30369)
OUTPUT(g34446)
OUTPUT(g29230)
OUTPUT(g34789)
OUTPUT(g3983)
OUTPUT(g33975)
OUTPUT(g30497)
OUTPUT(g31917)
OUTPUT(g30418)
OUTPUT(g25721)
OUTPUT(g34622)
OUTPUT(g30438)
OUTPUT(g34266)
OUTPUT(g30540)
OUTPUT(g6358)
OUTPUT(g32986)
OUTPUT(g25648)
OUTPUT(g33960)
OUTPUT(g34442)
OUTPUT(g4277)
OUTPUT(g30421)
OUTPUT(g33573)
OUTPUT(g34730)
OUTPUT(g24205)
OUTPUT(g4294)
OUTPUT(g6005)
OUTPUT(g1399)
OUTPUT(g32979)
OUTPUT(g25731)
OUTPUT(g28078)
OUTPUT(g34025)
OUTPUT(g25763)
OUTPUT(g30481)
OUTPUT(g1500)
OUTPUT(g31890)
OUTPUT(g30517)
OUTPUT(g30539)
OUTPUT(g34880)
OUTPUT(g24242)
OUTPUT(g30436)
OUTPUT(g29265)
OUTPUT(g32990)
OUTPUT(g24245)
OUTPUT(g25739)
OUTPUT(g30553)
OUTPUT(g26907)
OUTPUT(g24278)
OUTPUT(g26955)
OUTPUT(g24282)
OUTPUT(g29276)
OUTPUT(g31894)
OUTPUT(g33037)
OUTPUT(g26894)
OUTPUT(g25711)
OUTPUT(g34593)
OUTPUT(g25654)
OUTPUT(g33962)
OUTPUT(g34451)
OUTPUT(g34250)
OUTPUT(g5331)
OUTPUT(g29295)
OUTPUT(g26905)
OUTPUT(g25629)
OUTPUT(g34792)
OUTPUT(g5798)
OUTPUT(g25703)
OUTPUT(g4000)
OUTPUT(g32983)
OUTPUT(g3668)
OUTPUT(g30402)
OUTPUT(g25757)
OUTPUT(g1426)
OUTPUT(g4446)
OUTPUT(g33999)
OUTPUT(g24262)
OUTPUT(g25729)
OUTPUT(g6140)
OUTPUT(g30558)
OUTPUT(g34848)
OUTPUT(g881)
OUTPUT(g31892)
OUTPUT(g26901)
OUTPUT(g26961)
OUTPUT(g33039)
OUTPUT(g33059)
OUTPUT(g31899)
OUTPUT(g33007)
OUTPUT(g25720)
OUTPUT(g21891)
OUTPUT(g30462)
OUTPUT(g18422)
OUTPUT(g30487)
OUTPUT(g33058)
OUTPUT(g31916)
OUTPUT(g24261)
OUTPUT(g25730)
OUTPUT(g30531)
OUTPUT(g30506)
OUTPUT(g34804)
OUTPUT(g25747)
OUTPUT(g4005)
OUTPUT(g33601)
OUTPUT(g26922)
OUTPUT(g878)
OUTPUT(g25679)
OUTPUT(g29250)
OUTPUT(g30459)
OUTPUT(g1582)
OUTPUT(g33534)
OUTPUT(g30543)
OUTPUT(g29275)
OUTPUT(g34030)
OUTPUT(g34980)
OUTPUT(g30451)
OUTPUT(g25723)
OUTPUT(g25627)
OUTPUT(g34787)
OUTPUT(g4222)
OUTPUT(g30552)
OUTPUT(g34996)
OUTPUT(g30337)
OUTPUT(g24254)
OUTPUT(g24277)
OUTPUT(g29237)
OUTPUT(g30378)
OUTPUT(g31912)
OUTPUT(g25603)
OUTPUT(g33019)
OUTPUT(g33623)
OUTPUT(g25608)
OUTPUT(g29235)
OUTPUT(g31902)
OUTPUT(g29306)
OUTPUT(g28080)
OUTPUT(g33978)
OUTPUT(g26970)
OUTPUT(g25660)
OUTPUT(g25726)
OUTPUT(g29278)
OUTPUT(g34253)
OUTPUT(g29272)
OUTPUT(g33595)
OUTPUT(g33610)
OUTPUT(g33589)
OUTPUT(g34605)
OUTPUT(g30350)
OUTPUT(g25611)
OUTPUT(g26936)
OUTPUT(g33619)
OUTPUT(g3798)
OUTPUT(g34022)
OUTPUT(g34033)
OUTPUT(g34726)
OUTPUT(g31870)
OUTPUT(g33985)
OUTPUT(g29283)
OUTPUT(g34003)
OUTPUT(g5101)
OUTPUT(g25727)
OUTPUT(g25677)
OUTPUT(g34463)
OUTPUT(g33006)
OUTPUT(g29292)
OUTPUT(g30557)
OUTPUT(g33989)
OUTPUT(g28098)
OUTPUT(g33033)
OUTPUT(g3654)
OUTPUT(g34005)
OUTPUT(g26932)
OUTPUT(g30516)
OUTPUT(g33575)
OUTPUT(g33032)
OUTPUT(g6329)
OUTPUT(g31891)
OUTPUT(g30486)
OUTPUT(g34991)
OUTPUT(g25678)
OUTPUT(g30440)
OUTPUT(g4191)
OUTPUT(g1570)
OUTPUT(g26949)
OUTPUT(g30530)
OUTPUT(g30542)
OUTPUT(g4213)
OUTPUT(g25624)
OUTPUT(g30383)
OUTPUT(g33597)
OUTPUT(g34598)
OUTPUT(g26957)
OUTPUT(g26967)
OUTPUT(g3447)
OUTPUT(g28102)
OUTPUT(g30524)
OUTPUT(g25671)
OUTPUT(g26903)
OUTPUT(g30475)
OUTPUT(g34647)
OUTPUT(g30377)
OUTPUT(g33553)
OUTPUT(g21902)
OUTPUT(g31903)
OUTPUT(g25715)
OUTPUT(g33984)
OUTPUT(g33602)
OUTPUT(g28045)
OUTPUT(g34603)
OUTPUT(g33035)
OUTPUT(g4304)
OUTPUT(g24208)
OUTPUT(g1239)
OUTPUT(g34596)
OUTPUT(g28064)
OUTPUT(g34990)
OUTPUT(g24213)
OUTPUT(g31887)
OUTPUT(g33614)
OUTPUT(g31907)
OUTPUT(g33060)
OUTPUT(g30362)
OUTPUT(g31875)
OUTPUT(g33023)
OUTPUT(g25674)
OUTPUT(g26898)
OUTPUT(g25618)
OUTPUT(g30518)
OUTPUT(g28079)
OUTPUT(g6974)
OUTPUT(g3303)
OUTPUT(g26959)
OUTPUT(g34801)
OUTPUT(g26884)
OUTPUT(g25600)
OUTPUT(g26933)
OUTPUT(g28066)
OUTPUT(g33612)
OUTPUT(g5327)
OUTPUT(g24268)
OUTPUT(g25716)
OUTPUT(g25675)
OUTPUT(g26906)
OUTPUT(g24203)
OUTPUT(g24346)
OUTPUT(g24207)
OUTPUT(g25701)
OUTPUT(g29269)
OUTPUT(g34592)
OUTPUT(g28068)
OUTPUT(g34255)
OUTPUT(g30450)
OUTPUT(g30456)
OUTPUT(g32991)
OUTPUT(g6144)
OUTPUT(g24348)
OUTPUT(g34249)
OUTPUT(g25713)
OUTPUT(g31909)
OUTPUT(g30371)
OUTPUT(g29268)
OUTPUT(g29224)
OUTPUT(g859)
OUTPUT(g33017)
OUTPUT(g30339)
OUTPUT(g33967)
OUTPUT(g4194)
OUTPUT(g5276)
OUTPUT(g33559)
OUTPUT(g29255)
OUTPUT(g5452)
OUTPUT(g30368)
OUTPUT(g30375)
OUTPUT(g25732)
OUTPUT(g28052)
OUTPUT(g28089)
OUTPUT(g33055)
OUTPUT(g30392)
OUTPUT(g30343)
OUTPUT(g25657)
OUTPUT(g30523)
OUTPUT(g24233)
OUTPUT(g33018)
OUTPUT(g32976)
OUTPUT(g30349)
OUTPUT(g33067)
OUTPUT(g26900)
OUTPUT(g31883)
OUTPUT(g33034)
OUTPUT(g30551)
OUTPUT(g25667)
OUTPUT(g30452)
OUTPUT(g25612)
OUTPUT(g31874)
OUTPUT(g34719)
OUTPUT(g33607)
OUTPUT(g26923)
OUTPUT(g25746)
OUTPUT(g24211)
OUTPUT(g33050)
OUTPUT(g24341)
OUTPUT(g1056)
OUTPUT(g24201)
OUTPUT(g30463)
OUTPUT(g6486)
OUTPUT(g34464)
OUTPUT(g25710)
OUTPUT(g24243)
OUTPUT(g24335)
OUTPUT(g34611)
OUTPUT(g34262)
OUTPUT(g30546)
OUTPUT(g18527)
OUTPUT(g25591)
OUTPUT(g4414)
OUTPUT(g30347)
OUTPUT(g10384)
OUTPUT(g5283)
OUTPUT(g30556)
OUTPUT(g33020)
OUTPUT(g34589)
OUTPUT(g33562)
OUTPUT(g35002)
OUTPUT(g25610)
OUTPUT(g33015)
OUTPUT(g31896)
OUTPUT(g34004)
OUTPUT(g30428)
OUTPUT(g30485)
OUTPUT(g30422)
OUTPUT(g25606)
OUTPUT(g25714)
OUTPUT(g25680)
OUTPUT(g29294)
OUTPUT(g30423)
OUTPUT(g30529)
OUTPUT(g34028)
OUTPUT(g25724)
OUTPUT(g33587)
OUTPUT(g30460)
OUTPUT(g31910)
OUTPUT(g30401)
OUTPUT(g33990)
OUTPUT(g3976)
OUTPUT(g1075)
OUTPUT(g29309)
OUTPUT(g30411)
OUTPUT(g33546)
OUTPUT(g28085)
OUTPUT(g26904)
OUTPUT(g33556)
OUTPUT(g18093)
OUTPUT(g25722)
OUTPUT(g25605)
OUTPUT(g33062)
OUTPUT(g26893)
OUTPUT(g5313)
OUTPUT(g28050)
OUTPUT(g34626)
OUTPUT(g33583)
OUTPUT(g30472)
OUTPUT(g34454)
OUTPUT(g34850)
OUTPUT(g4019)
OUTPUT(g4537)
OUTPUT(g24272)
OUTPUT(g31906)
OUTPUT(g5681)
OUTPUT(g24214)
OUTPUT(g25718)
OUTPUT(g26909)
OUTPUT(g30406)
OUTPUT(g33569)
OUTPUT(g25694)
OUTPUT(g34628)
OUTPUT(g34458)
OUTPUT(g24240)
OUTPUT(g31918)
OUTPUT(g34634)
OUTPUT(g25700)
OUTPUT(g29293)
OUTPUT(g18421)
OUTPUT(g33009)
OUTPUT(g33603)
OUTPUT(g24355)
OUTPUT(g34268)
OUTPUT(g25691)
OUTPUT(g26890)
OUTPUT(g4449)
OUTPUT(g29264)
OUTPUT(g28072)
OUTPUT(g31900)
OUTPUT(g25712)
OUTPUT(g26956)
OUTPUT(g29271)
OUTPUT(g29304)
OUTPUT(g5654)
OUTPUT(g29261)
OUTPUT(g28063)
OUTPUT(g1116)
OUTPUT(g34027)
OUTPUT(g33961)
OUTPUT(g25672)
OUTPUT(g33604)
OUTPUT(g33025)
OUTPUT(g4207)
OUTPUT(g32995)
OUTPUT(g34624)
OUTPUT(g30415)
OUTPUT(g33536)
OUTPUT(g26888)
OUTPUT(g28055)
OUTPUT(g24238)
OUTPUT(g31921)
OUTPUT(g33600)
OUTPUT(g28105)
OUTPUT(g34721)
OUTPUT(g29307)
OUTPUT(g30345)
OUTPUT(g34453)
OUTPUT(g32980)
OUTPUT(g29238)
OUTPUT(g34639)
OUTPUT(g25695)
OUTPUT(g33057)
OUTPUT(g26969)
OUTPUT(g31879)
OUTPUT(g29253)
OUTPUT(g34021)
OUTPUT(g26895)
OUTPUT(g30413)
OUTPUT(g30549)
OUTPUT(g24347)
OUTPUT(g25758)
OUTPUT(g34808)
OUTPUT(g30501)
OUTPUT(g33969)
OUTPUT(g34440)
OUTPUT(g5969)
OUTPUT(g30433)
OUTPUT(g21900)
OUTPUT(g26921)
OUTPUT(g31893)
OUTPUT(g29270)
OUTPUT(g34878)
OUTPUT(g33038)
OUTPUT(g31865)
OUTPUT(g26926)
OUTPUT(g28083)
OUTPUT(g29209)
OUTPUT(g34797)
OUTPUT(g30478)
OUTPUT(g34724)
OUTPUT(g24212)
OUTPUT(g26883)
OUTPUT(g32985)
OUTPUT(g25761)
OUTPUT(g26886)
OUTPUT(g34796)
OUTPUT(g32982)
OUTPUT(g33561)
OUTPUT(g26880)
OUTPUT(g34591)
OUTPUT(g31884)
OUTPUT(g26931)
OUTPUT(g884)
OUTPUT(g5308)
OUTPUT(g34641)
OUTPUT(g34629)
OUTPUT(g33598)
OUTPUT(g33576)
OUTPUT(g34720)
OUTPUT(g26902)
OUTPUT(g29244)
OUTPUT(g30468)
OUTPUT(g26924)
OUTPUT(g25645)
OUTPUT(g33031)
OUTPUT(g29245)
OUTPUT(g29266)
OUTPUT(g30559)
OUTPUT(g6715)
OUTPUT(g34794)
OUTPUT(g28087)
OUTPUT(g5677)
OUTPUT(g30435)
OUTPUT(g3969)
OUTPUT(g25609)
OUTPUT(g28095)
OUTPUT(g28057)
OUTPUT(g34439)
OUTPUT(g34595)
OUTPUT(g1233)
OUTPUT(g34260)
OUTPUT(g33012)
OUTPUT(g32989)
OUTPUT(g34006)
OUTPUT(g34847)
OUTPUT(g5983)
OUTPUT(g365)
OUTPUT(g26910)
OUTPUT(g21722)
OUTPUT(g25658)
OUTPUT(g28043)
OUTPUT(g33021)
OUTPUT(g29251)
OUTPUT(g25665)
OUTPUT(g6697)
OUTPUT(g34456)
OUTPUT(g26968)
OUTPUT(g33991)
OUTPUT(g3443)
OUTPUT(g26930)
OUTPUT(g34599)
OUTPUT(g28082)
OUTPUT(g33557)
OUTPUT(g30511)
OUTPUT(g33045)
OUTPUT(g3096)
OUTPUT(g30379)
OUTPUT(g24267)
OUTPUT(g34020)
OUTPUT(g28100)
OUTPUT(g24249)
OUTPUT(g31908)
OUTPUT(g25592)
OUTPUT(g30382)
OUTPUT(g29285)
OUTPUT(g25644)
OUTPUT(g1227)
OUTPUT(g34992)
OUTPUT(g25662)
OUTPUT(g21896)
OUTPUT(g33563)
OUTPUT(g33622)
OUTPUT(g31876)
OUTPUT(g33582)
OUTPUT(g6711)
OUTPUT(g28086)
OUTPUT(g25744)
OUTPUT(g29262)
OUTPUT(g24270)
OUTPUT(g33581)
OUTPUT(g194)
OUTPUT(g26937)
OUTPUT(g34849)
OUTPUT(g28060)
OUTPUT(g33618)
OUTPUT(g34038)
OUTPUT(g6000)
OUTPUT(g34032)
OUTPUT(g31927)
OUTPUT(g31919)
OUTPUT(g34803)
OUTPUT(g34459)
OUTPUT(g30509)
OUTPUT(g34640)
OUTPUT(g3298)
OUTPUT(g28069)
OUTPUT(g21899)
OUTPUT(g31868)
OUTPUT(g26938)
OUTPUT(g25756)
OUTPUT(g30363)
OUTPUT(g30334)
OUTPUT(g33970)
OUTPUT(g30391)
OUTPUT(g25615)
OUTPUT(g33540)
OUTPUT(g30445)
OUTPUT(g25725)
OUTPUT(g25617)
OUTPUT(g24247)
OUTPUT(g24215)
OUTPUT(g3649)
OUTPUT(g33964)
OUTPUT(g25719)
OUTPUT(g29228)
OUTPUT(g30514)
OUTPUT(g33627)
OUTPUT(g28101)
OUTPUT(g24231)
OUTPUT(g34615)
OUTPUT(g30356)
OUTPUT(g25696)
OUTPUT(g30493)
OUTPUT(g4219)
OUTPUT(g33594)
OUTPUT(g34009)
OUTPUT(g30365)
OUTPUT(g33004)
OUTPUT(g34018)
OUTPUT(g25685)
OUTPUT(g34040)
OUTPUT(g25639)
OUTPUT(g34029)
OUTPUT(g30488)
OUTPUT(g34600)
OUTPUT(g29300)
OUTPUT(g6369)
OUTPUT(g34802)
OUTPUT(g25614)
OUTPUT(g28058)
OUTPUT(g29225)
OUTPUT(g33580)
OUTPUT(g30532)
OUTPUT(g6365)
OUTPUT(g5320)
OUTPUT(g25760)
OUTPUT(g25620)
OUTPUT(g4188)
OUTPUT(g33054)
OUTPUT(g26962)
OUTPUT(g33564)
OUTPUT(g32984)
OUTPUT(g34039)
OUTPUT(g31932)
OUTPUT(g33065)
OUTPUT(g30443)
OUTPUT(g29291)
OUTPUT(g24279)
OUTPUT(g30508)
OUTPUT(g29232)
OUTPUT(g34269)
OUTPUT(g30464)
OUTPUT(g33988)
OUTPUT(g30522)
OUTPUT(g25708)
OUTPUT(g5290)
OUTPUT(g30374)
OUTPUT(g26953)
OUTPUT(g34008)
OUTPUT(g34444)
OUTPUT(g34731)
OUTPUT(g33606)
OUTPUT(g24334)
OUTPUT(g34265)
OUTPUT(g30340)
OUTPUT(g24257)
OUTPUT(g30482)
OUTPUT(g25673)
OUTPUT(g31929)
OUTPUT(g34604)
OUTPUT(g3632)
OUTPUT(g33591)
OUTPUT(g4226)
OUTPUT(g30525)
OUTPUT(g26929)
OUTPUT(g30448)
OUTPUT(g34602)
OUTPUT(g30513)
OUTPUT(g30469)
OUTPUT(g33608)
OUTPUT(g33626)
OUTPUT(g34725)
OUTPUT(g30342)
OUTPUT(g29267)
OUTPUT(g25593)
OUTPUT(g30548)
OUTPUT(g33052)
OUTPUT(g34012)
OUTPUT(g34017)
OUTPUT(g34785)
OUTPUT(g24263)
OUTPUT(g26912)
OUTPUT(g30364)
OUTPUT(g34254)
OUTPUT(g34251)
OUTPUT(g30560)
OUTPUT(g33983)
OUTPUT(g25752)
OUTPUT(g6346)
OUTPUT(g6692)
OUTPUT(g24204)
OUTPUT(g33980)
OUTPUT(g34631)
OUTPUT(g28103)
OUTPUT(g31873)
OUTPUT(g29243)
OUTPUT(g25740)
OUTPUT(g25623)
OUTPUT(g26950)
OUTPUT(g4999)
OUTPUT(g30431)
OUTPUT(g30467)
OUTPUT(g30353)
OUTPUT(g34467)
OUTPUT(g30442)
OUTPUT(g29305)
OUTPUT(g25616)
OUTPUT(g29252)
OUTPUT(g1459)
OUTPUT(g6972)
OUTPUT(g4216)
OUTPUT(g33003)
OUTPUT(g34613)
OUTPUT(g4027)
OUTPUT(g33570)
OUTPUT(g4809)
OUTPUT(g33061)
OUTPUT(g21723)
OUTPUT(g34734)
OUTPUT(g24275)
OUTPUT(g4408)
OUTPUT(g887)
OUTPUT(g29302)
OUTPUT(g24349)
OUTPUT(g34264)
OUTPUT(g30484)
OUTPUT(g25634)
OUTPUT(g33567)
OUTPUT(g33585)
OUTPUT(g30527)
OUTPUT(g34995)
OUTPUT(g30447)
OUTPUT(g344)
OUTPUT(g31914)
OUTPUT(g34256)
OUTPUT(g25630)
OUTPUT(g29290)
OUTPUT(g29227)
OUTPUT(g31872)
OUTPUT(g29287)
OUTPUT(g31897)
OUTPUT(g6719)
OUTPUT(g30562)
OUTPUT(g34011)
OUTPUT(g33996)
OUTPUT(g21898)
OUTPUT(g33014)
OUTPUT(g34465)
OUTPUT(g33995)
OUTPUT(g30372)
OUTPUT(g30545)
OUTPUT(g30389)
OUTPUT(g33590)
OUTPUT(g34616)
OUTPUT(g26927)
OUTPUT(g32992)
OUTPUT(g3281)
OUTPUT(g25631)
OUTPUT(g30477)
OUTPUT(g34632)
OUTPUT(g28046)
OUTPUT(g4287)
OUTPUT(g26896)
OUTPUT(g25602)
OUTPUT(g26916)
OUTPUT(g33578)
OUTPUT(g25745)
OUTPUT(g4204)
OUTPUT(g33579)
OUTPUT(g30354)
OUTPUT(g30425)
OUTPUT(g24200)
OUTPUT(g33544)
OUTPUT(g25764)
OUTPUT(g31930)
OUTPUT(g24246)
OUTPUT(g30507)
OUTPUT(g26889)
OUTPUT(g30333)
OUTPUT(g215)
OUTPUT(g25753)
OUTPUT(g32998)
OUTPUT(g32987)
OUTPUT(g25702)
OUTPUT(g29286)
OUTPUT(g34606)
OUTPUT(g33070)
OUTPUT(g29240)
OUTPUT(g32999)
OUTPUT(g33605)
OUTPUT(g24255)
OUTPUT(g26945)
OUTPUT(g34877)
OUTPUT(g33558)
OUTPUT(g25647)
OUTPUT(g31889)
OUTPUT(g25699)
OUTPUT(g29289)
OUTPUT(g30388)
OUTPUT(g799)
OUTPUT(g29254)
OUTPUT(g28074)
OUTPUT(g34450)
OUTPUT(g30512)
OUTPUT(g33572)
OUTPUT(g5976)
OUTPUT(g15048)
OUTPUT(g33551)
OUTPUT(g33538)
OUTPUT(g33005)
OUTPUT(g24248)
OUTPUT(g33002)
OUTPUT(g24234)
OUTPUT(g30471)
OUTPUT(g34000)
OUTPUT(g34016)
OUTPUT(g33048)
OUTPUT(g26911)
OUTPUT(g5002)
OUTPUT(g18528)
OUTPUT(g6019)
OUTPUT(g25628)
OUTPUT(g26934)
OUTPUT(g31928)
OUTPUT(g869)
OUTPUT(g34468)
OUTPUT(g24202)
OUTPUT(g33542)
OUTPUT(g1422)
OUTPUT(g34717)
OUTPUT(g34445)
OUTPUT(g28104)
OUTPUT(g33555)
OUTPUT(g34013)
OUTPUT(g28091)
OUTPUT(g26919)
OUTPUT(g4812)
OUTPUT(g6322)
OUTPUT(g30554)
OUTPUT(g29281)
OUTPUT(g1079)
OUTPUT(g30537)
OUTPUT(g28092)
OUTPUT(g34732)
OUTPUT(g28049)
OUTPUT(g33545)
OUTPUT(g30441)
OUTPUT(g29247)
OUTPUT(g24354)
OUTPUT(g25636)
OUTPUT(g31911)
OUTPUT(g26914)
OUTPUT(g25670)
OUTPUT(g33998)
OUTPUT(g25626)
OUTPUT(g33977)
OUTPUT(g29297)
OUTPUT(g28071)
OUTPUT(g30387)
OUTPUT(g33577)
OUTPUT(g25737)
OUTPUT(g33592)
OUTPUT(g26913)
OUTPUT(g28044)
OUTPUT(g26948)
OUTPUT(g31931)
OUTPUT(g30344)
OUTPUT(g26885)
OUTPUT(g33069)
OUTPUT(g34621)
OUTPUT(g28075)
OUTPUT(g28059)
OUTPUT(g25762)
OUTPUT(g3274)
OUTPUT(g25646)
OUTPUT(g34633)
OUTPUT(g24352)
OUTPUT(g26925)
OUTPUT(g30446)
OUTPUT(g25597)
OUTPUT(g24342)
OUTPUT(g30357)
OUTPUT(g26908)
OUTPUT(g21905)
OUTPUT(g30399)
OUTPUT(g29242)
OUTPUT(g25659)
OUTPUT(g30547)
OUTPUT(g31881)
OUTPUT(g34010)
OUTPUT(g33986)
OUTPUT(g34257)
OUTPUT(g30544)
OUTPUT(g30561)
OUTPUT(g5005)
OUTPUT(g30430)
OUTPUT(g34799)
OUTPUT(g33565)
OUTPUT(g33968)
OUTPUT(g34879)
OUTPUT(g34793)
OUTPUT(g25754)
OUTPUT(g33566)
OUTPUT(g6661)
OUTPUT(g30465)
OUTPUT(g28073)
OUTPUT(g24351)
OUTPUT(g30346)
OUTPUT(g21893)
OUTPUT(g4815)
OUTPUT(g31904)
OUTPUT(g34635)
OUTPUT(g25637)
OUTPUT(g29274)
OUTPUT(g6675)
OUTPUT(g30396)
OUTPUT(g25735)
OUTPUT(g34037)
OUTPUT(g34791)
OUTPUT(g30520)
OUTPUT(g30358)
OUTPUT(g29299)
OUTPUT(g28081)
OUTPUT(g28096)
OUTPUT(g28088)
OUTPUT(g24241)
OUTPUT(g30397)
OUTPUT(g4520)
OUTPUT(g30409)
OUTPUT(g29284)
OUTPUT(g30470)
OUTPUT(g30367)
OUTPUT(g24273)
OUTPUT(g29288)
OUTPUT(g30359)
OUTPUT(g25698)
OUTPUT(g30398)
OUTPUT(g4023)
OUTPUT(g34718)
OUTPUT(g26952)
OUTPUT(g34590)
OUTPUT(g26928)
OUTPUT(g4197)
OUTPUT(g26954)
OUTPUT(g30351)
OUTPUT(g31871)
OUTPUT(g5105)
OUTPUT(g34594)
OUTPUT(g26939)
OUTPUT(g33994)
OUTPUT(g25596)
OUTPUT(g33586)
OUTPUT(g21901)
OUTPUT(g31866)
OUTPUT(g33000)
OUTPUT(g26918)
OUTPUT(g33051)
OUTPUT(g28065)
OUTPUT(g30373)
OUTPUT(g28056)
OUTPUT(g34601)
OUTPUT(g30355)
OUTPUT(g30426)
OUTPUT(g34805)
OUTPUT(g31913)
OUTPUT(g34002)
OUTPUT(g6704)
OUTPUT(g25652)
OUTPUT(g28053)
OUTPUT(g29229)
OUTPUT(g33620)
OUTPUT(g34722)
OUTPUT(g33599)
OUTPUT(g30515)
OUTPUT(g25649)
OUTPUT(g33066)
OUTPUT(g33979)
OUTPUT(g30417)
OUTPUT(g25683)
OUTPUT(g33574)
OUTPUT(g5673)
OUTPUT(g30410)
OUTPUT(g30454)
OUTPUT(g34024)
OUTPUT(g33547)
OUTPUT(g30386)
OUTPUT(g33596)
OUTPUT(g26887)
OUTPUT(g34607)
OUTPUT(g33056)
OUTPUT(g31895)
OUTPUT(g33068)
OUTPUT(g29233)
OUTPUT(g24258)
OUTPUT(g30376)
OUTPUT(g33549)
OUTPUT(g29308)
OUTPUT(g25759)
OUTPUT(g30408)
OUTPUT(g29241)
OUTPUT(g34620)
OUTPUT(g33621)
OUTPUT(g25707)
OUTPUT(g24339)
OUTPUT(g4185)
OUTPUT(g25738)
OUTPUT(g34443)
OUTPUT(g34619)
OUTPUT(g29234)
OUTPUT(g30503)
OUTPUT(g21724)
OUTPUT(g3310)
OUTPUT(g30550)
OUTPUT(g33001)
OUTPUT(g33040)
OUTPUT(g30492)
OUTPUT(g25664)
OUTPUT(g26944)
OUTPUT(g3672)
OUTPUT(g34614)
OUTPUT(g29260)
OUTPUT(g3325)
OUTPUT(g33047)
OUTPUT(g25692)
OUTPUT(g25733)
OUTPUT(g30536)
OUTPUT(g1157)
OUTPUT(g31888)
OUTPUT(g29246)
OUTPUT(g34261)
OUTPUT(g33611)
OUTPUT(g25638)
OUTPUT(g34728)
OUTPUT(g29222)
OUTPUT(g25742)
OUTPUT(g30449)
OUTPUT(g25643)
OUTPUT(g34608)
OUTPUT(g24345)
OUTPUT(g31922)
OUTPUT(g34994)
OUTPUT(g25635)
OUTPUT(g25686)
OUTPUT(g30461)
OUTPUT(g34466)
OUTPUT(g31901)
OUTPUT(g29249)
OUTPUT(g26882)
OUTPUT(g33041)
OUTPUT(g33011)
OUTPUT(g25734)
OUTPUT(g28097)
OUTPUT(g33030)
OUTPUT(g5659)
OUTPUT(g34618)
OUTPUT(g33010)
OUTPUT(g4229)
OUTPUT(g31864)
OUTPUT(g34630)
OUTPUT(g31898)
OUTPUT(g25653)
OUTPUT(g25632)
OUTPUT(g32988)
OUTPUT(g33616)
OUTPUT(g29280)
OUTPUT(g33609)
OUTPUT(g30563)
OUTPUT(g33044)
OUTPUT(g30437)
OUTPUT(g30412)
OUTPUT(g5630)
OUTPUT(g21725)
OUTPUT(g3267)
OUTPUT(g30491)
OUTPUT(g30434)
OUTPUT(g34612)
OUTPUT(g29259)
OUTPUT(g3321)
OUTPUT(g25681)
OUTPUT(g25687)
OUTPUT(g33617)
OUTPUT(g30479)
OUTPUT(g29256)
OUTPUT(g28054)
OUTPUT(g30535)
OUTPUT(g28094)
OUTPUT(g30385)
OUTPUT(g30361)
OUTPUT(g25705)
OUTPUT(g24260)
OUTPUT(g29257)
OUTPUT(g34461)
OUTPUT(g34258)
OUTPUT(g32993)
OUTPUT(g33992)
OUTPUT(g28061)
OUTPUT(g30394)
OUTPUT(g34449)
OUTPUT(g34019)
OUTPUT(g21726)
OUTPUT(g29231)
OUTPUT(g25682)
OUTPUT(g21897)
OUTPUT(g28067)
OUTPUT(g30395)
OUTPUT(g21892)
OUTPUT(g31885)
OUTPUT(g4210)
OUTPUT(g28048)
OUTPUT(g34723)
OUTPUT(g25717)
OUTPUT(g25598)
OUTPUT(g33987)
OUTPUT(g30380)
OUTPUT(g5448)
OUTPUT(g26965)
OUTPUT(g25706)
OUTPUT(g30458)
OUTPUT(g24338)
OUTPUT(g30400)
OUTPUT(g21904)
OUTPUT(g34623)
OUTPUT(g24343)
OUTPUT(g25666)
OUTPUT(g30473)
OUTPUT(g24252)
OUTPUT(g33028)
OUTPUT(g29258)
OUTPUT(g30407)
OUTPUT(g26958)
OUTPUT(g34457)
OUTPUT(g33568)
OUTPUT(g25663)
OUTPUT(g26964)
OUTPUT(g4200)
OUTPUT(g34735)
OUTPUT(g30352)
OUTPUT(g33543)
OUTPUT(g24271)
OUTPUT(g30326)
OUTPUT(g33981)
OUTPUT(g30500)
OUTPUT(g34786)
OUTPUT(g29277)
g9900(1) = NOT(g6)
g9954(3) = NAND(g6128, g6120)
g6895(4) = NOT(g3288)
g9797(2) = NOT(g5441)
g6837(1) = NOT(g968)
I15824(1) = NOT(g1116)
g10160(4) = NAND(g5623, g5666, g5637, g5659)
g9510(1) = NOT(g5835)
I13031(1) = NOT(g6747)
I12910(1) = NOT(g4340)
g10289(1) = NOT(g1319)
g7888(2) = NOT(g1536)
g9291(3) = NOT(g3021)
I13718(1) = NOT(g890)
g8224(2) = NOT(g3774)
I17932(1) = NOT(g3310)
I12530(1) = NOT(g4815)
g10308(2) = NOT(g4459)
g9902(1) = NOT(g100)
g9259(4) = NOT(g5176)
I15190(1) = NOT(g6005)
I12483(1) = NOT(g3096)
g9819(1) = NOT(g92)
g7297(3) = NOT(g6069)
I12779(1) = NOT(g4210)
g9488(1) = NOT(g1878)
g7138(1) = NOT(g5360)
g7963(1) = NOT(g4146)
g6903(1) = NOT(g3502)
g7109(1) = NOT(g5011)
I12199(1) = NOT(g6215)
g6854(1) = NOT(g2685)
g6941(4) = NOT(g3990)
g9951(2) = NOT(g6133)
I18600(1) = NOT(g5335)
g6989(1) = NOT(g4575)
g9152(1) = NOT(g2834)
g8945(2) = NOT(g608)
g7957(2) = NOT(g1252)
g7049(1) = NOT(g5853)
g6958(1) = NOT(g4372)
g7175(2) = NOR(g6098, g6058)
g8340(1) = NOT(g3050)
I12109(1) = NOT(g749)
g7715(1) = NOT(g1178)
g8478(1) = NOT(g3103)
g9594(1) = NOT(g2307)
g6829(1) = NOT(g1319)
g7498(1) = NOT(g6675)
g9806(1) = NOT(g5782)
I16741(1) = NOT(g5677)
I12855(1) = NOT(g4311)
g9887(1) = NOT(g5802)
I11746(1) = NOT(g4570)
g9934(1) = NOT(g5849)
g10042(1) = NOT(g2671)
I16803(1) = NOT(g6369)
I13321(1) = NOT(g6486)
I12884(1) = NOT(g4213)
I16391(1) = NOT(g859)
g7162(1) = NOT(g4521)
g7268(6) = NOT(g1636)
I11740(1) = NOT(g4519)
g7362(6) = NOT(g1906)
g9433(2) = NOT(g5148)
I13740(1) = NOT(g85)
I11685(1) = NOT(g117)
g8310(5) = NOT(g2051)
g6978(3) = NOT(g4616)
g9496(1) = NOT(g3303)
g8663(2) = NOT(g3343)
g10030(1) = NOT(g116)
I18614(1) = NOT(g6315)
g10093(2) = NOT(g5703)
g8107(4) = NOT(g3179)
g9891(2) = NOT(g6173)
g8002(2) = NOT(g1389)
g9337(1) = NOT(g1608)
g9913(1) = NOT(g2403)
g10185(4) = NAND(g5969, g6012, g5983, g6005)
g7086(1) = NOT(g4826)
g8236(1) = NOT(g4812)
g10108(1) = NOT(g120)
g10219(2) = NOT(g2697)
g9807(1) = NOT(g5712)
g6849(1) = NOT(g2551)
g10218(1) = NOT(g2527)
g7470(1) = NOT(g5623)
g10033(1) = NOT(g655)
g6900(2) = NOT(g3440)
g8928(4) = NOT(g4340)
g9815(1) = NOT(g6098)
g8064(3) = NOT(g3376)
g8899(3) = NOT(g807)
g8534(3) = NOT(g3338)
I11908(1) = NOT(g4449)
g9692(1) = NOT(g1756)
I12767(1) = NOT(g4197)
I13166(1) = NOT(g5101)
I12994(1) = NOT(g6748)
g9354(5) = NOT(g2719)
g9960(1) = NOT(g6474)
I16401(1) = NOT(g869)
g7635(1) = NOT(g1002)
I12189(1) = NOT(g5869)
g6819(1) = NOT(g1046)
g7087(4) = NOT(g6336)
g7487(2) = NOT(g1259)
g8237(1) = NOT(g255)
I18460(1) = NOT(g5276)
I12183(1) = NOT(g2719)
g6923(2) = NOT(g3791)
g10037(1) = NOT(g1848)
I12826(1) = NOT(g4349)
g9883(3) = NAND(g5782, g5774)
g6804(3) = NOT(g490)
g10155(1) = NOT(g2643)
g9761(1) = NOT(g2445)
g7192(2) = NOR(g6444, g6404)
I11992(1) = NOT(g763)
g6870(2) = NOT(g3089)
g9828(1) = NOT(g2024)
g8948(2) = NOT(g785)
g6825(1) = NOT(g979)
g7369(4) = NOT(g1996)
g8955(1) = NOT(g1418)
g10194(2) = NOT(g6741)
I18504(1) = NOT(g5283)
g8356(1) = NOT(g54)
I16371(1) = NOT(g887)
g7868(1) = NOT(g1099)
I15102(1) = NOT(g5313)
I11835(1) = NOT(g101)
I13326(1) = NOT(g66)
g8150(3) = NOT(g2185)
g7041(4) = NOT(g5644)
g8350(2) = NOT(g4646)
g7535(1) = NOT(g1500)
I13007(1) = NOT(g65)
I12360(1) = NOT(g528)
g10119(1) = NOT(g2841)
g8438(1) = NOT(g3100)
g8009(1) = NOT(g3106)
g7261(1) = NOT(g4449)
g10118(1) = NOT(g2541)
g9932(1) = NOT(g5805)
I16829(1) = NOT(g6715)
g8836(2) = NOT(g736)
g6887(1) = NOT(g3333)
I12893(1) = NOT(g4226)
g7246(1) = NOT(g4446)
g10053(3) = NOT(g6381)
g9576(4) = NOT(g6565)
g8229(4) = NOT(g3881)
g9716(4) = NOT(g5057)
g8993(4) = NOT(g385)
g10036(1) = NOT(g1816)
g8822(6) = NOT(g4975)
g10177(1) = NOT(g1834)
I13684(1) = NOT(g128)
g9848(3) = NOT(g4462)
I19837(1) = NOT(g1399)
g6845(1) = NOT(g2126)
g9699(1) = NOT(g2311)
I13329(1) = NOT(g86)
g9766(4) = NOT(g2748)
I15717(1) = NOT(g6346)
g10074(3) = NOT(g718)
I12159(1) = NOT(g608)
g7216(2) = NOT(g822)
I11785(1) = NOT(g5703)
g8895(2) = NOT(g599)
g10166(2) = NOT(g6040)
g9644(1) = NOT(g2016)
g8620(2) = NOT(g3065)
g8462(3) = NOT(g1183)
g7247(3) = NOT(g5377)
I12046(1) = NOT(g613)
g7564(1) = NOT(g336)
I18509(1) = NOT(g5623)
g9818(1) = NOT(g6490)
g6815(1) = NOT(g929)
I12787(1) = NOT(g4311)
I12776(1) = NOT(g4207)
g8249(5) = NOT(g1917)
I15238(1) = NOT(g6351)
I13010(1) = NOT(g6749)
g6960(1) = NOT(g1)
g9386(3) = NOT(g5727)
I18813(1) = NOT(g5673)
g7308(5) = NOT(g1668)
I12382(1) = NOT(g47)
g9599(1) = NOT(g3310)
g9274(5) = NOT(g5857)
g9614(1) = NOT(g5128)
I18647(1) = NOT(g5320)
g9543(2) = NAND(g2217, g2185)
g8854(3) = NOT(g613)
g9821(1) = NOT(g115)
I13236(1) = NOT(g5452)
I16168(1) = NOT(g3321)
I17857(1) = NOT(g3969)
I13054(1) = NOT(g6744)
g9326(5) = NOT(g6203)
g10176(1) = NOT(g44)
I16217(1) = NOT(g3632)
g9311(4) = NOT(g5523)
g10154(2) = NOT(g2547)
g9083(2) = NOT(g626)
I16639(1) = NOT(g4000)
g8219(4) = NOT(g3731)
g9636(1) = NOT(g72)
g7827(1) = NOT(g4688)
g9705(2) = NAND(g2619, g2587)
g8431(2) = NOT(g3085)
I15663(1) = NOT(g5308)
I12805(1) = NOT(g4098)
g6828(1) = NOT(g1300)
I18333(1) = NOT(g1083)
I12890(1) = NOT(g4219)
g8632(2) = NAND(g1514, g1500)
g6830(1) = NOT(g1389)
g8005(3) = NOT(g3025)
I11860(1) = NOT(g43)
g7582(3) = NAND(g1361, g1373)
I12572(1) = NOT(g51)
g9187(6) = NOT(g518)
I15677(1) = NOT(g5654)
I12003(1) = NOT(g767)
g8286(1) = NOT(g53)
g8765(1) = NOT(g3333)
g7780(1) = NOT(g2878)
g8912(1) = NOT(g4180)
g9200(2) = NOT(g1548)
g8733(1) = NOT(g3698)
g7018(4) = NOT(g5297)
I12930(1) = NOT(g4349)
I11726(1) = NOT(g4273)
g7418(4) = NOT(g2361)
I13726(1) = NOT(g4537)
g9003(3) = NOT(g790)
g6953(1) = NOT(g4157)
I12336(1) = NOT(g52)
g8125(4) = NOT(g3869)
g6956(1) = NOT(g4242)
g8796(6) = NOT(g4785)
g10083(1) = NOT(g2407)
g8324(5) = NOT(g2476)
I16417(1) = NOT(g875)
I13252(1) = NOT(g6751)
g8540(1) = NOT(g3408)
g9223(2) = NOT(g1216)
g7197(3) = NOT(g812)
I16762(1) = NOT(g5290)
g6848(1) = NOT(g2417)
g7397(3) = NOT(g890)
g10139(1) = NOT(g136)
g6855(1) = NOT(g2711)
g8287(2) = NOT(g160)
g9416(1) = NOT(g2429)
I13037(1) = NOT(g4304)
I11635(1) = NOT(g9)
g8399(1) = NOT(g3798)
g8728(4) = NAND(g3618, g3661, g3632, g3654)
I12026(1) = NOT(g344)
g8898(1) = NOT(g676)
g7631(1) = NOT(g74)
I11903(1) = NOT(g4414)
g7301(2) = NOT(g925)
I12503(1) = NOT(g215)
g6818(1) = NOT(g976)
g9880(2) = NOT(g5787)
I12523(1) = NOT(g3794)
g9537(1) = NOT(g1748)
g7751(1) = NOT(g1521)
g8259(7) = NOT(g2217)
g10200(2) = NOT(g2138)
g9978(3) = NOT(g2756)
I12811(1) = NOT(g4340)
g10115(1) = NOT(g2283)
I18662(1) = NOT(g6322)
g8088(2) = NOT(g1554)
g6975(1) = NOT(g4507)
I13124(1) = NOT(g2729)
g7964(5) = NOT(g3155)
I13483(1) = NOT(g6035)
I13606(1) = NOT(g74)
g7441(1) = NOT(g862)
g9982(1) = NOT(g3976)
g9234(4) = NOT(g5170)
I11750(1) = NOT(g4474)
I12451(1) = NOT(g3092)
g9542(1) = NOT(g2173)
I11655(1) = NOT(g1246)
g8951(2) = NOT(g554)
g6984(1) = NOT(g4709)
I17814(1) = NOT(g3274)
g8114(4) = NOT(g3522)
g10184(1) = NOT(g4486)
I18778(1) = NOT(g6704)
g9554(1) = NOT(g5105)
I12837(1) = NOT(g4222)
g8650(1) = NOT(g4664)
I12896(1) = NOT(g4229)
I13020(1) = NOT(g6750)
g7411(6) = NOT(g2040)
g8136(1) = NOT(g269)
g8594(1) = NOT(g3849)
I11623(1) = NOT(g28)
I11801(1) = NOT(g6395)
g7002(1) = NOT(g5160)
I11980(1) = NOT(g66)
g7992(1) = NOT(g5008)
g9490(1) = NOT(g2563)
I14563(1) = NOT(g802)
g9166(7) = NOT(g837)
g6904(1) = NOT(g3494)
I12112(1) = NOT(g794)
g9056(3) = NOT(g3017)
g9456(3) = NOT(g6073)
g8228(1) = NOT(g3835)
g9529(4) = NOT(g6561)
g7863(3) = NOT(g1249)
g9800(3) = NAND(g5436, g5428)
I12997(1) = NOT(g351)
I14395(1) = NOT(g3654)
g6841(3) = NOT(g2145)
g8033(3) = NOT(g157)
g9698(1) = NOT(g2181)
g9964(1) = NOT(g126)
g9591(2) = NAND(g1926, g1894)
I12793(1) = NOT(g4578)
g8195(5) = NOT(g1783)
g8137(1) = NOT(g411)
g8891(3) = NOT(g582)
I16193(1) = NOT(g3281)
g7266(1) = NOT(g35)
g9595(2) = NAND(g2351, g2319)
g8807(1) = NOT(g79)
g9619(1) = NOT(g5845)
g7400(3) = NOT(g911)
g8859(3) = NOT(g772)
g6811(2) = NOT(g714)
g7601(9) = NOR(g1322, g1333)
g7092(2) = NOT(g6483)
I13634(1) = NOT(g79)
g9843(4) = NOT(g4311)
g9989(2) = NOT(g5077)
g7063(1) = NOT(g4831)
g6874(1) = NOT(g3143)
I12519(1) = NOT(g3447)
g9834(1) = NOT(g2579)
g9971(1) = NOT(g2093)
g9686(1) = NOT(g73)
g8255(3) = NOT(g2028)
g7183(1) = NOT(g4608)
I12618(1) = NOT(g3338)
I12128(1) = NOT(g4253)
g9598(1) = NOT(g2571)
g8097(4) = NOT(g3029)
g7779(1) = NOT(g1413)
g8497(2) = NOT(g3436)
g8154(2) = NOT(g3139)
g8354(1) = NOT(g4815)
g7023(2) = NOT(g5445)
g10206(1) = NOT(g4489)
g9321(4) = NOT(g5863)
g7423(1) = NOT(g2433)
g9670(1) = NOT(g5022)
g7846(3) = NAND(g4843, g4878)
I11843(1) = NOT(g111)
g7361(1) = NOT(g1874)
g10114(1) = NOT(g2116)
g9253(3) = NOT(g5037)
I16821(1) = NOT(g5983)
g10082(1) = NOT(g2375)
I11793(1) = NOT(g6049)
g9909(1) = NOT(g1978)
I12761(1) = NOT(g4188)
g7451(4) = NOT(g2070)
g6982(1) = NOT(g4531)
g7327(1) = NOT(g2165)
g8112(1) = NOT(g3419)
g8218(2) = NOT(g3490)
g9740(1) = NOT(g5821)
g8267(5) = NOT(g2342)
I18276(1) = NOT(g1075)
I12120(1) = NOT(g632)
g9552(1) = NOT(g3654)
g7017(1) = NOT(g128)
I11820(1) = NOT(g3869)
g8676(1) = NOT(g4821)
g6999(2) = NOT(g86)
g6800(1) = NOT(g203)
I13152(1) = NOT(g6746)
I13287(1) = NOT(g110)
I18752(1) = NOT(g6358)
g8830(2) = NOT(g767)
g8592(1) = NOT(g3805)
g7072(1) = NOT(g6199)
I11691(1) = NOT(g36)
g7472(1) = NOT(g6329)
g9860(1) = NOT(g5417)
g7046(2) = NOT(g5791)
g7443(2) = NOT(g914)
I12709(1) = NOT(g4284)
g7116(1) = NOT(g22)
I13875(1) = NOT(g1233)
g9691(2) = NOT(g1706)
I12056(1) = NOT(g2748)
g8068(1) = NOT(g3457)
g9607(5) = NOT(g5046)
g9962(2) = NOT(g6519)
g9158(3) = NOT(g513)
g8677(1) = NOT(g4854)
g7533(1) = NOT(g1306)
g9506(2) = NOT(g5774)
I18555(1) = NOT(g5630)
g7697(3) = NOT(g4087)
I12070(1) = NOT(g785)
I13708(1) = NOT(g136)
g10106(1) = NOT(g16)
I11743(1) = NOT(g4564)
I12887(1) = NOT(g4216)
g8848(3) = NOT(g358)
I15208(1) = NOT(g637)
I12563(1) = NOT(g3798)
g9444(4) = NOT(g5535)
g9174(2) = NOT(g1205)
I18835(1) = NOT(g6365)
g9374(4) = NOT(g5188)
I15542(1) = NOT(g1570)
g6918(4) = NOT(g3639)
g7936(2) = NOT(g1061)
g9985(3) = NOT(g4332)
g9856(3) = NOT(g5343)
I12764(1) = NOT(g4194)
g8241(7) = NOT(g1792)
I11816(1) = NOT(g93)
I12132(1) = NOT(g577)
g9284(1) = NOT(g2161)
g7202(6) = NOT(g4639)
g9239(5) = NOT(g5511)
g9180(3) = NOT(g3719)
g9380(1) = NOT(g5471)
g9832(2) = NOT(g2399)
g10109(1) = NOT(g135)
I16575(1) = NOT(g3298)
g9853(2) = NOT(g5297)
g8644(2) = NOT(g3352)
g9020(2) = NOT(g4287)
g7922(3) = NOT(g1312)
g8119(3) = NOT(g3727)
g10338(2) = NOR(g5062, g5022)
g8751(4) = NAND(g3969, g4012, g3983, g4005)
g8571(1) = NOT(g57)
g7581(1) = NOT(g1379)
g9559(4) = NOT(g6077)
I11737(1) = NOT(g4467)
I12808(1) = NOT(g4322)
g9931(1) = NOT(g5763)
g7597(1) = NOT(g952)
g7611(3) = NAND(g4057, g4064)
I16606(1) = NOT(g3649)
g8211(3) = NOT(g2319)
g9905(1) = NOT(g802)
g9407(5) = NOT(g6549)
g8186(1) = NOT(g990)
I13552(1) = NOT(g121)
g9630(1) = NOT(g6527)
g7995(2) = NOT(g153)
g8026(5) = NOT(g3857)
g7479(7) = NOT(g1008)
g9300(4) = NOT(g5180)
g8426(4) = NOT(g3045)
g8170(1) = NOT(g3770)
g7840(1) = NOT(g4878)
g6827(1) = NOT(g1277)
I16875(1) = NOT(g6675)
g10121(1) = NOT(g2327)
g8280(1) = NOT(g3443)
g9973(1) = NOT(g2112)
g7356(4) = NOT(g1802)
I17819(1) = NOT(g3618)
g9040(3) = NOT(g499)
I13672(1) = NOT(g106)
g9969(1) = NOT(g1682)
I18845(1) = NOT(g6711)
I12167(1) = NOT(g5176)
g8106(1) = NOT(g3133)
g8187(7) = NOT(g1657)
g8387(1) = NOT(g3080)
g7163(2) = NOT(g4593)
I13548(1) = NOT(g94)
g8756(1) = NOT(g4049)
g9648(1) = NOT(g2177)
g10028(1) = NOT(g8)
g9875(4) = NOT(g5747)
I12086(1) = NOT(g622)
g8046(5) = NOT(g528)
g8514(1) = NOT(g4258)
g7985(5) = NOT(g3506)
I12568(1) = NOT(g5005)
g8345(1) = NOT(g3794)
I12823(1) = NOT(g4311)
g7157(1) = NOT(g5706)
I12749(1) = NOT(g4575)
g9839(2) = NOT(g2724)
I13723(1) = NOT(g3167)
I13149(1) = NOT(g6745)
I16847(1) = NOT(g6329)
I11620(1) = NOT(g1)
I12144(1) = NOT(g554)
I18709(1) = NOT(g6668)
g9618(1) = NOT(g5794)
g8858(1) = NOT(g671)
g9282(1) = NOT(g723)
g8016(4) = NOT(g3391)
I12746(1) = NOT(g4087)
I12580(1) = NOT(g1239)
g9693(1) = NOT(g1886)
g6985(1) = NOT(g4669)
I12631(1) = NOT(g1242)
g8522(3) = NOT(g298)
I13206(1) = NOT(g5448)
I15536(1) = NOT(g1227)
g6995(1) = NOT(g4944)
g9804(1) = NOT(g5456)
g10262(3) = NOT(g586)
g10224(4) = NAND(g6661, g6704, g6675, g6697)
g9792(4) = NOT(g5401)
I11665(1) = NOT(g1589)
g7778(1) = NOT(g1339)
g8654(1) = NOT(g1087)
g9621(4) = NOT(g6423)
g10191(2) = NOT(g6386)
I11896(1) = NOT(g4446)
I18337(1) = NOT(g1422)
I12861(1) = NOT(g4372)
I12666(1) = NOT(g4040)
I11716(1) = NOT(g4054)
g7475(3) = NOT(g896)
g7627(3) = NOT(g4311)
I11708(1) = NOT(g3703)
g8612(3) = NOT(g2775)
g9518(4) = NOT(g6219)
I12013(1) = NOT(g590)
g7998(3) = NOT(g392)
g6986(1) = NOT(g4743)
I18728(1) = NOT(g6012)
g9776(1) = NOT(g5073)
g10099(2) = NOT(g6682)
I12954(1) = NOT(g4358)
g6983(1) = NOT(g4698)
g7439(1) = NOT(g6351)
g8130(1) = NOT(g4515)
I12644(1) = NOT(g3689)
g8330(3) = NOT(g2587)
I13705(1) = NOT(g63)
g9965(1) = NOT(g127)
g9264(4) = NOT(g5396)
g9360(3) = NOT(g3372)
g9933(1) = NOT(g5759)
g10032(1) = NOT(g562)
g10140(1) = NOT(g19)
g9050(1) = NOT(g1087)
g7952(1) = NOT(g3774)
g9450(1) = NOT(g5817)
I14450(1) = NOT(g4191)
I12016(1) = NOT(g772)
I13581(1) = NOT(g6727)
I11777(1) = NOT(g5357)
g9379(1) = NOT(g5424)
g6836(1) = NOT(g1322)
I18700(1) = NOT(g6027)
I11697(1) = NOT(g3352)
g9777(1) = NOT(g5112)
g7503(7) = NOT(g1351)
g7970(1) = NOT(g4688)
g8056(1) = NOT(g1246)
I13317(1) = NOT(g6144)
g8456(1) = NOT(g56)
I16357(1) = NOT(g884)
g8155(4) = NOT(g3380)
g7224(2) = NOT(g4601)
I12534(1) = NOT(g50)
g8851(2) = NOT(g590)
I13057(1) = NOT(g112)
g6839(1) = NOT(g1858)
g8964(2) = NOT(g4269)
I11626(1) = NOT(g31)
g9100(2) = NOR(g3752, g3712)
g9569(4) = NOT(g6227)
I12030(1) = NOT(g595)
g9541(1) = NOT(g2012)
I12089(1) = NOT(g744)
g9332(1) = NOT(g64)
I13276(1) = NOT(g5798)
I12991(1) = NOT(g6752)
g10147(3) = NOT(g728)
g6816(1) = NOT(g933)
I12487(1) = NOT(g3443)
g9744(1) = NOT(g6486)
g7095(1) = NOT(g6545)
g6988(1) = NOT(g4765)
g9748(1) = NOT(g114)
g8872(1) = NOT(g4258)
g10151(1) = NOT(g1992)
g10172(2) = NOT(g6459)
g7892(4) = NOT(g4801)
g9558(2) = NOT(g5841)
g8057(1) = NOT(g3068)
g8744(1) = NOT(g691)
g8457(1) = NOT(g225)
I12935(1) = NOT(g6753)
g6994(1) = NOT(g4933)
g9901(1) = NOT(g84)
I12927(1) = NOT(g4332)
g9511(4) = NOT(g5881)
I12176(1) = NOT(g5523)
g8686(3) = NOT(g2819)
g7991(1) = NOT(g4878)
g7244(1) = NOT(g4408)
g9492(4) = NOT(g2759)
g7340(2) = NOT(g4443)
g9600(1) = NOT(g3632)
g9574(1) = NOT(g6462)
I13424(1) = NOT(g5689)
g7907(1) = NOT(g3072)
g8626(3) = NOT(g4040)
g9714(1) = NOT(g4012)
g10059(1) = NOT(g6451)
g7517(1) = NOT(g962)
g9392(4) = NOT(g5869)
g10058(1) = NOT(g6497)
g7876(2) = NOT(g1495)
g8938(5) = NOT(g4899)
g10203(1) = NOT(g2393)
I16181(1) = NOT(g3672)
g10044(2) = NOT(g5357)
g8519(2) = NOT(g287)
I12735(1) = NOT(g4572)
I12418(1) = NOT(g55)
g6940(1) = NOT(g4035)
g8606(1) = NOT(g4653)
g10120(1) = NOT(g1902)
I11753(1) = NOT(g4492)
g9889(1) = NOT(g6128)
g7110(4) = NOT(g6682)
g10072(1) = NOT(g9)
g7824(2) = NOT(g4169)
g6996(1) = NOT(g4955)
g9602(4) = NOR(g4688, g4681, g4674, g4646)
g7236(2) = NOT(g4608)
g9285(5) = NOT(g2715)
g9500(2) = NOT(g5495)
g8341(1) = NOT(g3119)
g7549(3) = NAND(g1018, g1030)
g9184(1) = NOT(g6120)
g9339(1) = NOT(g2295)
g9024(5) = NOT(g4358)
g7040(1) = NOT(g4821)
g7222(1) = NOT(g4427)
g9809(5) = NOT(g6082)
g9581(1) = NOT(g91)
I18825(1) = NOT(g6019)
g7928(3) = NOT(g4776)
I12858(1) = NOT(g4340)
g8607(1) = NOT(g37)
g9664(4) = NOR(g4878, g4871, g4864, g4836)
g7064(4) = NOT(g5990)
g9672(5) = NOT(g5390)
g9077(5) = NOT(g504)
g8659(3) = NOT(g2815)
I12541(1) = NOT(g194)
g8506(1) = NOT(g3782)
g9523(3) = NOT(g6419)
g7785(2) = NOT(g4621)
I17964(1) = NOT(g3661)
g6799(1) = NOT(g199)
g8587(3) = NOT(g3689)
g9689(1) = NOT(g124)
g7948(3) = AND(g1548, g1430)
g7563(1) = NOT(g6322)
g6997(1) = NOT(g4578)
g9551(1) = NOT(g3281)
g9742(1) = NOT(g6144)
I12987(1) = NOT(g12)
g9099(1) = NOT(g3706)
g9499(1) = NOT(g5152)
I12064(1) = NOT(g617)
g7394(1) = NOT(g5637)
g9051(3) = NOT(g1426)
g8434(3) = NAND(g3080, g3072)
g9654(2) = NAND(g2485, g2453)
I14619(1) = NOT(g4185)
g9754(1) = NOT(g2020)
g6802(1) = NOT(g468)
g8284(1) = NOT(g5002)
g8239(1) = NOT(g1056)
g10181(1) = NOT(g2551)
g7557(1) = NOT(g1500)
g8180(1) = NOT(g262)
g8591(1) = NOT(g3763)
g9613(1) = NOT(g5062)
g7471(1) = NOT(g6012)
g9044(3) = NOT(g604)
g9269(4) = NOT(g5517)
g8507(1) = NOT(g3712)
g9983(1) = NOT(g4239)
g9862(1) = NOT(g5413)
g7139(2) = NOR(g5406, g5366)
g10190(1) = NOT(g6044)
g9206(5) = NOT(g5164)
g9724(3) = NAND(g5092, g5084)
I12712(1) = NOT(g59)
I12907(1) = NOT(g4322)
g9534(1) = NOT(g90)
g9729(1) = NOT(g5138)
g9961(1) = NOT(g6404)
g7438(1) = NOT(g5983)
g8630(1) = NOT(g4843)
g9927(3) = NOT(g5689)
g8300(1) = NOT(g1242)
I18667(1) = NOT(g6661)
g9014(1) = NOT(g3004)
g10102(3) = NOT(g6727)
g9414(1) = NOT(g2004)
g7212(3) = NOT(g6411)
g9660(1) = NOT(g3267)
g9946(4) = NOT(g6093)
g9903(1) = NOT(g681)
I12092(1) = NOT(g790)
I12333(1) = NOT(g45)
g10274(1) = NOT(g976)
g9036(1) = NOT(g5084)
g8440(1) = NOT(g3431)
g9679(1) = NOT(g5475)
g8123(1) = NOT(g3808)
g9831(1) = NOT(g2269)
g8666(2) = NOT(g3703)
g10060(1) = NOT(g6541)
g10197(1) = NOT(g31)
g9805(1) = NOT(g5485)
g9916(1) = NOT(g3625)
I13892(1) = NOT(g1576)
I12577(1) = NOT(g1227)
g9749(1) = NOT(g1691)
I18560(1) = NOT(g5969)
g8655(3) = NOT(g2787)
g7462(6) = NOT(g2599)
g6838(1) = NOT(g1724)
g6809(1) = NOT(g341)
I12083(1) = NOT(g568)
I12819(1) = NOT(g4277)
g7788(2) = NOT(g4674)
g9095(3) = NOT(g3368)
g9037(2) = NOT(g164)
g9653(1) = NOT(g2441)
g8172(4) = NOT(g3873)
g8278(1) = NOT(g3096)
g10111(1) = NOT(g1858)
g9995(3) = NOT(g6035)
g7392(1) = NOT(g4438)
I12463(1) = NOT(g4812)
g8343(1) = NOT(g3447)
g9752(2) = NOT(g1840)
g8282(2) = NOT(g3841)
g8566(1) = NOT(g3831)
I13473(1) = NOT(g4157)
g7854(2) = NOT(g1152)
I12415(1) = NOT(g48)
I13374(1) = NOT(g6490)
g8334(5) = NOT(g3034)
g6926(1) = NOT(g3853)
I11617(1) = NOT(g1)
g8804(1) = NOT(g4035)
g10150(1) = NOT(g1700)
g9364(4) = NOT(g5041)
I12963(1) = NOT(g640)
I12790(1) = NOT(g4340)
g7219(2) = NOT(g4405)
g10019(2) = NOT(g6479)
g7431(4) = NOT(g2555)
g7252(4) = NOT(g1592)
I12214(1) = NOT(g6561)
g8113(1) = NOT(g3466)
I18092(1) = NOT(g3668)
g7405(4) = NOT(g1936)
I13202(1) = NOT(g5105)
g7765(1) = NOT(g4165)
I12608(1) = NOT(g1582)
I11734(1) = NOT(g4473)
g8567(3) = NOT(g4082)
g7733(4) = NOT(g4093)
I15697(1) = NOT(g6000)
g6927(1) = NOT(g3845)
g10001(1) = NOT(g6105)
g9888(1) = NOT(g5831)
g10077(1) = NOT(g1724)
g8593(1) = NOT(g3759)
g7073(1) = NOT(g6191)
I12799(1) = NOT(g59)
g9429(3) = NOT(g3723)
g7473(1) = NOT(g6697)
I16713(1) = NOT(g5331)
I11721(1) = NOT(g4145)
g7980(4) = NOT(g3161)
g7069(2) = NOT(g6137)
I15284(1) = NOT(g6697)
g8160(2) = NOT(g3423)
g10157(1) = NOT(g2036)
g8450(1) = NOT(g3821)
g9684(1) = NOT(g6191)
g8967(3) = NAND(g4264, g4258)
g9745(1) = NOT(g6537)
g9639(1) = NOT(g1752)
g9338(1) = NOT(g1870)
g10231(1) = NOT(g2661)
g9963(1) = NOT(g7)
g6831(1) = NOT(g1413)
g9309(1) = NOT(g5462)
g8179(1) = NOT(g4999)
g9808(2) = NOT(g5827)
g9759(2) = NOT(g2265)
g7898(4) = NOT(g4991)
I18653(1) = NOT(g5681)
I12538(1) = NOT(g58)
g9049(1) = NOT(g640)
g9449(1) = NOT(g5770)
g8609(2) = NAND(g1171, g1157)
g9575(1) = NOT(g6509)
g8165(4) = NOT(g3530)
g7344(1) = NOT(g5659)
g9498(1) = NOT(g5101)
g6873(1) = NOT(g3151)
g9833(1) = NOT(g2449)
I13715(1) = NOT(g71)
g7259(1) = NOT(g4375)
g8997(2) = NOT(g577)
g10085(1) = NOT(g1768)
g8541(1) = NOT(g3498)
I12411(1) = NOT(g4809)
g8680(1) = NOT(g686)
I13623(1) = NOT(g4294)
g6917(1) = NOT(g3684)
g9162(3) = NOT(g622)
I12950(1) = NOT(g4287)
I18609(1) = NOT(g5976)
g7886(1) = NOT(g1442)
I13352(1) = NOT(g4146)
g10156(1) = NOT(g2675)
g8558(2) = NOT(g3787)
g7314(1) = NOT(g1740)
g10180(1) = NOT(g2259)
g10175(1) = NOT(g28)
g7870(2) = NOT(g1193)
g10335(1) = NOT(g4483)
g7650(4) = NOT(g4064)
I18360(1) = NOT(g1426)
g8561(3) = NAND(g3782, g3774)
g9086(4) = NOT(g847)
g9728(1) = NOT(g5109)
g9730(1) = NOT(g5436)
g8092(1) = NOT(g1589)
I16795(1) = NOT(g5637)
g8492(4) = NOT(g3396)
g9070(1) = NOT(g5428)
g8714(1) = NOT(g4859)
g7972(2) = NOT(g1046)
g7806(2) = NOT(g4681)
g7943(2) = NOT(g1395)
I12758(1) = NOT(g4093)
g7322(4) = NOT(g1862)
g6990(1) = NOT(g4742)
g10278(2) = NOT(g4628)
I11701(1) = NOT(g4164)
g9678(1) = NOT(g5406)
g10039(1) = NOT(g2273)
g8623(2) = NOT(g3990)
I11809(1) = NOT(g6741)
g10038(1) = NOT(g2241)
I12141(1) = NOT(g599)
I13280(1) = NOT(g6140)
g7096(1) = NOT(g6537)
g9305(3) = NOT(g5381)
g7496(1) = NOT(g5969)
g7845(1) = NOT(g1146)
g7195(1) = NOT(g25)
g7395(1) = NOT(g6005)
g7891(1) = NOT(g2994)
g8651(2) = NOT(g758)
g7913(2) = NOT(g1052)
I12135(1) = NOT(g807)
g10143(3) = NOT(g568)
I12497(1) = NOT(g49)
g9226(2) = NOT(g1564)
I17787(1) = NOT(g3267)
g10169(2) = NOT(g6395)
g6808(1) = NOT(g554)
g8139(6) = NOT(g1648)
I12049(1) = NOT(g781)
g9373(1) = NOT(g5142)
g9091(1) = NOT(g1430)
g9491(1) = NOT(g2729)
g9822(1) = NOT(g125)
g10217(1) = NOT(g2102)
g9283(1) = NOT(g1736)
g9369(2) = NOT(g5084)
g9007(3) = NOT(g1083)
g6957(1) = NOT(g2932)
I11892(1) = NOT(g4408)
g8672(1) = NOT(g4669)
g9920(3) = NOT(g4322)
I15144(1) = NOT(g5659)
g8477(1) = NOT(g3061)
g7497(1) = NOT(g6358)
g9582(2) = NOT(g703)
g7960(2) = NOT(g1404)
g8205(5) = NOT(g2208)
g10223(1) = NOT(g4561)
I12106(1) = NOT(g626)
I12605(1) = NOT(g1570)
g8364(1) = NOT(g1585)
g8742(1) = NOT(g4035)
I16246(1) = NOT(g3983)
g10084(1) = NOT(g2837)
g9415(1) = NOT(g2169)
g10110(1) = NOT(g661)
I12033(1) = NOT(g776)
g7267(1) = NOT(g1604)
g10178(1) = NOT(g2126)
g9721(2) = NOT(g5097)
g8273(3) = NOT(g2453)
g7293(2) = NOT(g4452)
I18758(1) = NOT(g6719)
I17999(1) = NOT(g4012)
I18107(1) = NOT(g4019)
I13637(1) = NOT(g102)
g7828(2) = NOT(g4871)
I12654(1) = NOT(g1585)
g10334(1) = NOT(g4420)
g7592(1) = NOT(g347)
g9671(2) = NOT(g5134)
g9030(5) = NOT(g4793)
g9247(2) = NOT(g1559)
g7953(3) = NOT(g4966)
g9564(2) = NOT(g6120)
g9826(1) = NOT(g1844)
g10117(1) = NOT(g2509)
g10000(1) = NOT(g6151)
g8903(1) = NOT(g1075)
g9910(2) = NOT(g2108)
g9638(1) = NOT(g1620)
g7716(1) = NOT(g1199)
g7149(1) = NOT(g4564)
g7349(2) = NOT(g1270)
I12437(1) = NOT(g4999)
g6801(1) = NOT(g391)
I17938(1) = NOT(g3676)
g10124(4) = NAND(g5276, g5320, g5290, g5313)
I13694(1) = NOT(g117)
g9861(1) = NOT(g5459)
g10318(1) = NOR(g25, g22)
g8691(4) = NAND(g3267, g3310, g3281, g3303)
g9827(2) = NOT(g1974)
g9333(2) = NOT(g417)
I15036(1) = NOT(g799)
I16201(1) = NOT(g4023)
g7258(1) = NOT(g4414)
g7577(3) = NOT(g1263)
g7867(1) = NOT(g1489)
g9061(2) = NOR(g3401, g3361)
g10014(4) = NOT(g6439)
g10073(1) = NOT(g134)
I18795(1) = NOT(g5327)
I12172(1) = NOT(g2715)
I11688(1) = NOT(g70)
g8292(3) = NAND(g218, g215)
g8037(1) = NOT(g405)
I13360(1) = NOT(g5343)
g8102(2) = NOT(g3072)
g8302(7) = NOT(g1926)
I18297(1) = NOT(g1418)
g8579(3) = NOT(g2771)
g7975(4) = NOT(g3040)
g10116(2) = NOT(g2413)
g9662(1) = NOT(g3983)
g9018(1) = NOT(g4273)
I12719(1) = NOT(g365)
g7026(1) = NOT(g5507)
g9467(4) = NOT(g6434)
I12770(1) = NOT(g4200)
I15837(1) = NOT(g1459)
g7170(3) = NOT(g5719)
g10275(2) = NOT(g4584)
g9816(1) = NOT(g6167)
g7280(4) = NOT(g2153)
g7939(3) = NOT(g1280)
g8442(2) = NOT(g3476)
g10035(2) = NOT(g1720)
I12899(1) = NOT(g4232)
g7544(3) = NOT(g918)
g8164(1) = NOT(g3484)
g9381(4) = NOT(g5527)
g7636(3) = NOT(g4098)
g9685(2) = NOT(g6533)
g9197(2) = NOT(g1221)
g9397(4) = NOT(g6088)
g8770(3) = NOT(g749)
g8296(1) = NOT(g246)
g8725(2) = NOT(g739)
g7187(3) = NOT(g6065)
g7387(4) = NOT(g2421)
g7461(1) = NOT(g2567)
g8553(4) = NOT(g3747)
g10130(2) = NOT(g5694)
g6850(3) = NOT(g2704)
g7027(1) = NOT(g5499)
I19818(1) = NOT(g1056)
g10165(1) = NOT(g5698)
I18694(1) = NOT(g5666)
g9631(4) = NOT(g6573)
g8389(2) = NOT(g3125)
g7446(3) = NOT(g1256)
g7514(1) = NOT(g6704)
I14424(1) = NOT(g4005)
g8990(2) = NOT(g146)
g9257(1) = NOT(g5115)
g7003(1) = NOT(g5152)
I13539(1) = NOT(g6381)
g8171(1) = NOT(g3817)
g7345(3) = NOT(g6415)
g7841(3) = NOT(g904)
I12773(1) = NOT(g4204)
g6826(1) = NOT(g218)
g10222(1) = NOT(g4492)
g7191(1) = NOT(g6398)
g9751(1) = NOT(g1710)
g8281(1) = NOT(g3494)
g7536(1) = NOT(g5976)
g9585(1) = NOT(g1616)
g8297(2) = NOT(g142)
g7858(4) = NOT(g947)
I12061(1) = NOT(g562)
g8745(2) = NOT(g744)
g8138(1) = NOT(g1500)
g8639(3) = NOT(g2807)
g9645(2) = NAND(g2060, g2028)
g7522(1) = NOT(g6661)
g7115(1) = NOT(g12)
g8808(3) = NOT(g595)
g7315(6) = NOT(g1772)
g9669(1) = NOT(g5092)
I17852(1) = NOT(g3625)
g7158(2) = NOR(g5752, g5712)
g8201(3) = NOT(g1894)
g9890(1) = NOT(g6058)
g8449(1) = NOT(g3752)
g9011(1) = NOT(g1422)
g6846(1) = NOT(g2152)
g8575(3) = NOT(g291)
g7880(4) = NOT(g1291)
g8715(2) = NOT(g4927)
I12067(1) = NOT(g739)
g6803(1) = NOT(g496)
g7537(2) = NOT(g311)
g8833(2) = NOT(g794)
g9992(2) = NOT(g5990)
g8584(2) = NOT(g3639)
g8539(1) = NOT(g3454)
g9863(1) = NOT(g5503)
I12355(1) = NOT(g46)
g9480(2) = NOT(g559)
g9713(1) = NOT(g3618)
g10320(2) = NOT(g817)
g7328(6) = NOT(g2197)
g8362(1) = NOT(g194)
I13744(1) = NOT(g3518)
I12151(1) = NOT(g604)
g8052(2) = NOT(g1211)
g9688(1) = NOT(g113)
g6847(1) = NOT(g2283)
g9976(1) = NOT(g2537)
g10153(1) = NOT(g2417)
g8504(1) = NOT(g3451)
g10136(2) = NOT(g6113)
g9000(2) = NOT(g632)
I12227(1) = NOT(g34)
g8070(4) = NOT(g3518)
g7512(1) = NOT(g5283)
g9760(1) = NOT(g2315)
g7490(4) = NOT(g2629)
g9071(1) = NOT(g2831)
g7166(1) = NOT(g4311)
g7456(4) = NOT(g2495)
g6817(1) = NOT(g956)
g7649(1) = NOT(g1345)
g9924(2) = NOT(g5644)
g9220(2) = NOT(g843)
g7851(2) = NOT(g921)
g9779(1) = NOT(g5156)
g8406(1) = NOT(g232)
g8635(3) = NOT(g2783)
g9977(2) = NOT(g2667)
g8766(2) = NOT(g572)
g8087(1) = NOT(g1157)
g8748(2) = NOT(g776)
g9451(4) = NOT(g5873)
g9999(1) = NOT(g6109)
g7118(2) = NOT(g832)
g7619(1) = NOT(g1296)
g9103(1) = NOT(g5774)
I17892(1) = NOT(g3325)
I14365(1) = NOT(g3303)
g8373(7) = NOT(g2485)
g8091(2) = NOT(g1579)
I11629(1) = NOT(g19)
g7393(1) = NOT(g5320)
g6987(1) = NOT(g4754)
g9732(2) = NOT(g5481)
g9753(1) = NOT(g1890)
I12493(1) = NOT(g5002)
g7971(1) = NOT(g4818)
g7686(2) = NOT(g4659)
g8407(3) = NOT(g1171)
g9072(1) = NOT(g2994)
g8059(4) = NOT(g3171)
g9472(4) = NOT(g6555)
I11682(1) = NOT(g2756)
g8718(1) = NOT(g3333)
g9443(1) = NOT(g5489)
g7670(3) = NOT(g4104)
g9316(4) = NOT(g5742)
g6992(1) = NOT(g4899)
g9434(4) = NOT(g5385)
g7232(2) = NOT(g4411)
g7909(3) = NOT(g936)
I12103(1) = NOT(g572)
I18734(1) = NOT(g6373)
g9681(1) = NOT(g5798)
g10040(1) = NOT(g2652)
g7519(1) = NOT(g1157)
g9914(2) = NOT(g2533)
g7567(9) = NOR(g979, g990)
g9820(1) = NOT(g99)
g9462(4) = NOT(g6215)
g9413(1) = NOT(g1744)
g10183(1) = NOT(g2595)
I16770(1) = NOT(g6023)
g8388(1) = NOT(g3010)
g8216(1) = NOT(g3092)
g9601(1) = NOT(g4005)
I16328(1) = NOT(g878)
g10213(2) = NOT(g6732)
g9060(1) = NOT(g3355)
g9460(1) = NOT(g6154)
I15732(1) = NOT(g6692)
g8741(1) = NOT(g4821)
g10047(2) = NOT(g5421)
g10311(1) = NOT(g4633)
g9739(1) = NOT(g5752)
I13240(1) = NOT(g5794)
g7275(4) = NOT(g1728)
g8883(5) = NOT(g4709)
g7174(1) = NOT(g6052)
I17970(1) = NOT(g4027)
g7374(4) = NOT(g2227)
g8217(1) = NOT(g3143)
g9390(1) = NOT(g5808)
g8466(3) = NOT(g1514)
g9501(4) = NOT(g5731)
g7239(3) = NOT(g5033)
g8365(7) = NOT(g2060)
g7380(6) = NOT(g2331)
g10152(2) = NOT(g2122)
g7591(1) = NOT(g6668)
g8055(2) = NOT(g1236)
g9704(1) = NOT(g2575)
g8133(1) = NOT(g4809)
g8774(3) = NOT(g781)
g8396(1) = NOT(g3401)
g9250(1) = NOT(g1600)
g8538(1) = NOT(g3412)
I18066(1) = NOT(g3317)
g8509(4) = NOT(g4141)
I17901(1) = NOT(g3976)
I12000(1) = NOT(g582)
g9568(1) = NOT(g6181)
I16345(1) = NOT(g881)
g8418(7) = NOT(g2619)
g8290(1) = NOT(g218)
g9485(2) = NAND(g1657, g1624)
g8093(3) = NOT(g1624)
g10113(1) = NOT(g2084)
g7750(1) = NOT(g1070)
g8181(1) = NOT(g424)
g8381(5) = NOT(g2610)
g8685(1) = NOT(g1430)
g7440(1) = NOT(g329)
g8700(2) = NOT(g4054)
g8397(1) = NOT(g3470)
g9626(2) = NOT(g6466)
g8021(4) = NOT(g3512)
g6820(1) = NOT(g1070)
g7666(3) = NOT(g4076)
g7528(3) = NOT(g930)
g9683(1) = NOT(g6140)
g7655(3) = NOT(g4332)
g9778(1) = NOT(g5069)
g8631(1) = NOT(g283)
g10027(1) = NOT(g6523)
g8301(1) = NOT(g1399)
g7410(1) = NOT(g2008)
g9661(1) = NOT(g3661)
I12300(1) = NOT(g1157)
g10204(1) = NOT(g2685)
g10081(2) = NOT(g2279)
g8441(1) = NOT(g3361)
g7235(1) = NOT(g4521)
g7343(1) = NOT(g5290)
g9484(1) = NOT(g1612)
g9439(2) = NOT(g5428)
g6840(1) = NOT(g1992)
g8673(2) = NOT(g4737)
g7693(2) = NOT(g4849)
g7134(3) = NOT(g5029)
g7548(1) = NOT(g1036)
g8669(2) = NOT(g3767)
g10090(2) = NOT(g5348)
I13699(1) = NOT(g4581)
g10182(2) = NOT(g2681)
g8058(1) = NOT(g3115)
g8531(2) = NOT(g3288)
g8458(2) = NOT(g294)
g8743(1) = NOT(g550)
g8890(2) = NOT(g376)
g8505(1) = NOT(g3480)
g9616(1) = NOT(g5452)
g8011(4) = NOT(g3167)
g8734(2) = NOT(g4045)
g6954(1) = NOT(g4138)
g6810(1) = NOT(g723)
g9527(1) = NOT(g6500)
I12314(1) = NOT(g1500)
g7908(1) = NOT(g4157)
g8500(3) = NAND(g3431, g3423)
g10026(1) = NOT(g6494)
g9546(1) = NOT(g2437)
g10212(1) = NOT(g6390)
g7518(1) = NOT(g1024)
g9970(1) = NOT(g1714)
g8080(4) = NOT(g3863)
g8480(1) = NOT(g3147)
g8713(1) = NOT(g4826)
g7933(2) = NOT(g907)
g7521(1) = NOT(g5630)
g7050(1) = NOT(g5845)
g9516(1) = NOT(g6116)
g7231(1) = NOT(g5)
g9771(1) = NOT(g3969)
g9299(1) = NOT(g5124)
g9547(3) = NOT(g2735)
g7379(1) = NOT(g2299)
g8400(2) = NOT(g4836)
g9892(5) = NOT(g6428)
I11632(1) = NOT(g16)
g7289(3) = NOT(g4382)
g10133(2) = NOT(g6049)
g7835(1) = NOT(g4125)
g10229(1) = NOT(g6736)
I18293(1) = NOT(g1079)
g9015(2) = NOR(g3050, g3010)
g8806(1) = NAND(g358, g370, g376, g385)
g8183(2) = NOT(g482)
g8608(1) = NOT(g278)
I13094(1) = NOT(g2724)
g9907(1) = NOT(g1959)
g9959(1) = NOT(g6177)
g8977(6) = NOT(g4349)
g9517(1) = NOT(g6163)
g9690(1) = NOT(g732)
g7541(1) = NOT(g344)
g6998(1) = NOT(g4932)
g10112(2) = NOT(g1988)
g7132(1) = NOT(g4558)
g10050(2) = NOT(g6336)
g7153(3) = NOT(g5373)
g7680(4) = NOT(g4108)
g8451(4) = NOT(g4057)
g7701(2) = NAND(g4859, g4849, g4843)
g9915(1) = NOT(g2583)
g7802(1) = NOT(g324)
g8146(3) = NOT(g1760)
g10096(2) = NOT(g5767)
g8346(1) = NOT(g3845)
g9214(2) = NOT(g617)
I12041(1) = NOT(g2741)
g8696(1) = NOT(g3347)
g10207(4) = NAND(g6315, g6358, g6329, g6351)
g8508(2) = NOT(g3827)
g9402(4) = NOT(g6209)
g9824(1) = NOT(g1825)
g8944(1) = NOT(g370)
g8240(1) = NOT(g1333)
g8443(5) = NOT(g3736)
g9590(1) = NOT(g1882)
g9657(3) = NOT(g2763)
g8316(7) = NOT(g2351)
g9556(1) = NOT(g5448)
g8565(1) = NOT(g3802)
g10129(1) = NOT(g5352)
g9064(5) = NOT(g4983)
g8681(3) = NOT(g763)
g10002(1) = NOT(g6195)
g10057(1) = NOT(g6455)
g9899(1) = NOT(g6513)
g7262(3) = NOT(g5723)
g8697(2) = NOT(g3694)
g8914(1) = NOT(g4264)
g9194(2) = NOT(g827)
g10232(1) = NOT(g4527)
g7285(3) = NOT(g4643)
g9731(1) = NOT(g5366)
g9489(1) = NOT(g2303)
g9557(1) = NOT(g5499)
g10261(1) = NOT(g4555)
g7424(6) = NOT(g2465)
g7809(2) = NOT(g4864)
I12117(1) = NOT(g586)
g6991(1) = NOT(g4888)
g7523(2) = NOT(g305)
g7643(3) = NOT(g4322)
g9538(2) = NAND(g1792, g1760)
g6959(1) = NOT(g4420)
I12123(1) = NOT(g758)
g8479(1) = NOT(g3057)
g10080(1) = NOT(g1982)
g8840(2) = NOT(g4277)
g9212(1) = NOT(g6466)
g8390(5) = NOT(g3385)
g7926(1) = NOT(g3423)
g9229(4) = NOT(g5052)
g10199(1) = NOT(g1968)
g7918(3) = AND(g1205, g1087)
g10022(3) = NAND(g6474, g6466)
g8954(1) = NOT(g1079)
g8363(1) = NOT(g239)
g7534(1) = NOT(g1367)
g9620(2) = NOT(g6187)
g7927(1) = NOT(g4064)
g7836(3) = NAND(g4653, g4688)
I13597(1) = NOT(g4417)
g7903(3) = NOT(g969)
g10043(1) = NOT(g1632)
g7513(1) = NOT(g6315)
g9842(1) = NOT(g3274)
g9298(1) = NOT(g5080)
g7178(4) = NOT(g4392)
g7436(1) = NOT(g5276)
g7335(4) = NOT(g2287)
g7690(2) = NAND(g4669, g4659, g4653)
g10337(1) = NOT(g5016)
g7805(1) = NOT(g4366)
g7749(1) = NOT(g996)
g9708(4) = NOT(g2741)
g7947(1) = NOT(g1500)
g9252(2) = NOT(g4304)
g9958(1) = NOT(g6148)
g8075(4) = NOT(g3742)
g9829(1) = NOT(g2250)
g6814(1) = NOT(g632)
g7873(2) = NOT(g1266)
g10079(1) = NOT(g1950)
g9911(1) = NOT(g2384)
g7495(1) = NOT(g4375)
g7437(1) = NOT(g5666)
g10078(2) = NOT(g1854)
g8526(3) = NOT(g1526)
g9733(5) = NOT(g5736)
g10086(1) = NOT(g2193)
g9974(1) = NOT(g2518)
g7752(1) = NOT(g1542)
g8439(1) = NOT(g3129)
g9073(3) = NOT(g150)
g7917(1) = NOT(g1157)
g10159(1) = NOT(g4477)
g10158(1) = NOT(g2461)
g6993(1) = NOT(g4859)
g7932(1) = OR(g4072, g4153)
g7296(1) = NOT(g5313)
g8616(3) = NOT(g2803)
g7532(1) = NOT(g1157)
g7553(3) = NOT(g1274)
g8404(1) = NOT(g5005)
g8647(2) = NOT(g3416)
g8764(1) = NOT(g4826)
g9898(1) = NOT(g6444)
g8690(1) = AND(g2941, g2936)
g7764(1) = OR(g2999, g2932)
g8679(1) = OR(g222, g199)
g8720(1) = NOR(g358, g365)
g7396(1) = AND(g392, g441)
g10290(4) = AND(g4358, g4349)
g7685(1) = AND(g4382, g4375)
g8769(1) = NAND(g691, g714)
g7696(1) = AND(g2955, g2950)
g7834(1) = OR(g2886, g2946)
g8234(1) = AND(g4515, g4521)
g9984(1) = OR(g4300, g4242)
g9968(1) = AND(g1339, g1500)
g7499(2) = NOR(g333, g355)
g7684(1) = OR(g4072, g4176)
g7450(1) = OR(g1277, g1283)
g8530(1) = AND(g2902, g2907)
g7520(1) = AND(g2704, g2697, g2689)
g10123(1) = NOR(g4294, g4297)
g7469(1) = AND(g4382, g4438)
g8933(4) = NOR(g4709, g4785)
g7404(1) = OR(g933, g939)
g9535(1) = OR(g209, g538)
g8643(1) = AND(g2927, g2922)
g8984(4) = NOR(g4899, g4975)
g9217(2) = AND(g632, g626)
g8721(4) = AND(g385, g376, g365)
g7850(1) = NAND(g554, g807)
g7763(1) = AND(g2965, g2960)
g7251(1) = AND(g452, g392)
g8182(1) = NOR(g405, g392)
g10034(1) = AND(g1521, g1500)
g8461(1) = OR(g301, g534)
g9479(1) = AND(g305, g324)
g7804(1) = AND(g2975, g2970)
g9906(1) = AND(g996, g1157)
g7777(1) = AND(g723, g822, g817)
g7511(1) = AND(g2145, g2138, g2130)
g7781(3) = NOR(g4064, g4057)
g9967(1) = AND(g1178, g1157)
g7673(1) = OR(g4153, g4172)
g8583(1) = AND(g2917, g2912)
I12902(1) = OR(g4235, g4232, g4229, g4226)
I12903(1) = OR(g4222, g4219, g4216, g4213)
I12583(1) = OR(g1157, g1239, g990)
g9483(1) = OR(g1008, g969)
g9536(1) = OR(g1351, g1312)
I12611(1) = OR(g1500, g1582, g1333)
I12782(1) = OR(g4188, g4194, g4197, g4200)
I12783(1) = OR(g4204, g4207, g4210, g4180)
g8904(1) = OR(g1779, g1798)
g8905(1) = OR(g2204, g2223)
g9012(1) = OR(g2047, g2066)
g9055(1) = OR(g2606, g2625)
g8956(1) = OR(g1913, g1932)
g8957(1) = OR(g2338, g2357)
g9013(1) = OR(g2472, g2491)
g8863(1) = OR(g1644, g1664)
I13442(2) = NAND(g262, g239)
I12344(2) = NAND(g3106, g3111)
g9852(1) = NAND(g3684, g4871)
g9694(3) = NOR(g1936, g1862)
g9334(2) = NAND(g827, g832)
g7142(5) = NOR(g6573, g6565)
I13109(2) = NAND(g5808, g5813)
g7352(3) = NOR(g1526, g1514)
I12840(2) = NAND(g4222, g4235)
g9640(3) = NOR(g1802, g1728)
g8678(2) = NAND(g376, g358)
I13334(2) = NAND(g1687, g1691)
g8958(5) = NOR(g3881, g3873)
I12251(2) = NAND(g1124, g1129)
g10266(5) = NOR(g5188, g5180)
g10341(5) = NOR(g6227, g6219)
I13749(2) = NAND(g4608, g4584)
I13390(2) = NAND(g1821, g1825)
I13509(2) = NAND(g2089, g2093)
g8177(1) = NOR(g4966, g4991, g4983)
I12203(2) = NAND(g1094, g1135)
g9755(3) = NOR(g2070, g1996)
g7227(1) = NAND(g4584, g4593)
g9762(3) = NOR(g2495, g2421)
g8906(5) = NOR(g3530, g3522)
g8829(1) = NAND(g5011, g4836)
g7661(4) = NOR(g1211, g1216, g1221, g1205)
I13452(2) = NAND(g1955, g1959)
I13564(2) = NAND(g2648, g2652)
I13462(2) = NAND(g2380, g2384)
I12096(2) = NAND(g1339, g1322)
g9629(1) = NAND(g6462, g6466)
I12848(2) = NAND(g4281, g4277)
g8847(1) = NAND(g4831, g4681)
g8803(1) = NAND(g128, g4646)
g7228(2) = NAND(g6398, g6444)
g10281(5) = NOR(g5535, g5527)
g7150(2) = NAND(g5016, g5062)
I12728(2) = NAND(g4291, g4287)
I13182(2) = NAND(g6500, g6505)
g8105(1) = NAND(g3068, g3072)
I12261(2) = NAND(g1454, g1448)
I13729(2) = NAND(g4534, g4537)
I12269(2) = NAND(g1141, g956)
g7675(4) = NOR(g1554, g1559, g1564, g1548)
g9649(3) = NOR(g2227, g2153)
g9177(2) = NAND(g3355, g3401)
g9700(3) = NOR(g2361, g2287)
g9586(3) = NOR(g1668, g1592)
I12876(2) = NAND(g4200, g4180)
I11824(2) = NAND(g4593, g4601)
I12544(2) = NAND(g191, g194)
g9835(3) = NOR(g2629, g2555)
g9372(1) = NAND(g5080, g5084)
g8864(5) = NOR(g3179, g3171)
I12287(2) = NAND(g1484, g1300)
g9567(1) = NAND(g6116, g6120)
I12372(2) = NAND(g3457, g3462)
g10312(5) = NOR(g5881, g5873)
I12217(2) = NAND(g1437, g1478)
I12468(2) = NAND(g405, g392)
g9092(2) = NAND(g3004, g3050)
I12277(2) = NAND(g1467, g1472)
I13497(2) = NAND(g255, g232)
I12074(2) = NAND(g996, g979)
I12401(2) = NAND(g3808, g3813)
g8163(1) = NAND(g3419, g3423)
I13043(2) = NAND(g5115, g5120)
I11877(2) = NAND(g4388, g4430)
g7442(1) = NAND(g896, g890)
I13077(2) = NAND(g5462, g5467)
g9442(1) = NAND(g5424, g5428)
I11864(2) = NAND(g4434, g4401)
I13382(2) = NAND(g269, g246)
I13065(2) = NAND(g4308, g4304)
g9715(1) = NAND(g5011, g4836)
I12240(2) = NAND(g1111, g1105)
g9775(1) = NAND(g4831, g4681)
g9663(1) = NAND(g128, g4646)
I13401(2) = NAND(g2246, g2250)
g9246(1) = NAND(g847, g812)
g8889(1) = NAND(g3684, g4871)
g7167(2) = NAND(g5360, g5406)
g9203(2) = NAND(g3706, g3752)
I13518(2) = NAND(g2514, g2518)
g7304(3) = NOR(g1183, g1171)
g9509(1) = NAND(g5770, g5774)
g8227(1) = NAND(g3770, g3774)
I13139(2) = NAND(g6154, g6159)
g7184(2) = NAND(g5706, g5752)
g7209(2) = NAND(g6052, g6098)
g8131(1) = NOR(g4776, g4801, g4793)
g8347(2) = NAND(g4358, g4349, g4340)
g8086(1) = NOR(g168, g174, g182)
g10179(1) = NOR(g2098, g1964, g1830, g1696)
g10205(1) = NOR(g2657, g2523, g2389, g2255)
g7243(1) = NOT(I11892)
g7245(1) = NOT(I11896)
g7257(1) = NOT(I11903)
g7260(1) = NOT(I11908)
g7540(1) = NOT(I12026)
g7916(1) = NOT(I12300)
g7946(1) = NOT(I12314)
g8132(1) = NOT(I12411)
g8178(1) = NOT(I12437)
g8215(1) = NOT(I12451)
g8235(1) = NOT(I12463)
g8277(1) = NOT(I12483)
g8279(1) = NOT(I12487)
g8283(1) = NOT(I12493)
g8291(1) = NOT(I12503)
g8342(1) = NOT(I12519)
g8344(1) = NOT(I12523)
g8353(1) = NOT(I12530)
g8358(1) = NOT(I12541)
g8398(1) = NOT(I12563)
g8403(1) = NOT(I12568)
g8416(1) = NOT(I12580)
g8475(1) = NOT(I12608)
g8719(1) = NOT(I12719)
g8783(1) = NOT(I12761)
g8784(1) = NOT(I12764)
g8785(1) = NOT(I12767)
g8786(1) = NOT(I12770)
g8787(1) = NOT(I12773)
g8788(1) = NOT(I12776)
g8789(1) = NOT(I12779)
g8839(1) = NOT(I12819)
g8870(1) = NOT(I12837)
g8915(1) = NOT(I12884)
g8916(1) = NOT(I12887)
g8917(1) = NOT(I12890)
g8918(1) = NOT(I12893)
g8919(1) = NOT(I12896)
g8920(1) = NOT(I12899)
g9019(1) = NOT(I12950)
g9048(1) = NOT(I12963)
g9251(1) = NOT(I13037)
g9497(1) = NOT(I13166)
g9553(1) = NOT(I13202)
g9555(1) = NOT(I13206)
g9615(1) = NOT(I13236)
g9617(1) = NOT(I13240)
g9680(1) = NOT(I13276)
g9682(1) = NOT(I13280)
g9741(1) = NOT(I13317)
g9743(1) = NOT(I13321)
g9817(1) = NOT(I13374)
g10122(1) = NOT(I13623)
g10306(1) = NOT(I13726)
g10500(1) = NOT(I13875)
g10527(1) = NOT(I13892)
g11349(1) = NOT(I14365)
g11388(1) = NOT(I14395)
g11418(1) = NOT(I14424)
g11447(1) = NOT(I14450)
g11678(1) = NOT(I14563)
g11770(1) = NOT(I14619)
g12184(1) = NOT(I15036)
g12238(1) = NOT(I15102)
g12300(1) = NOT(I15144)
g12350(1) = NOT(I15190)
g12368(1) = NOT(I15208)
g12422(1) = NOT(I15238)
g12470(1) = NOT(I15284)
g12919(1) = NOT(I15536)
g12923(1) = NOT(I15542)
g13039(1) = NOT(I15663)
g13049(1) = NOT(I15677)
g13068(1) = NOT(I15697)
g13085(1) = NOT(I15717)
g13099(1) = NOT(I15732)
g13259(1) = NOT(I15824)
g13272(1) = NOT(I15837)
g13865(1) = NOT(I16168)
g13881(1) = NOT(I16181)
g13895(1) = NOT(I16193)
g13906(1) = NOT(I16201)
g13926(1) = NOT(I16217)
g13966(1) = NOT(I16246)
g14096(1) = NOT(I16328)
g14125(1) = NOT(I16345)
g14147(1) = NOT(I16357)
g14167(1) = NOT(I16371)
g14189(1) = NOT(I16391)
g14201(1) = NOT(I16401)
g14217(1) = NOT(I16417)
g14421(1) = NOT(I16575)
g14451(1) = NOT(I16606)
g14518(1) = NOT(I16639)
g14597(1) = NOT(I16713)
g14635(1) = NOT(I16741)
g14662(1) = NOT(I16762)
g14673(1) = NOT(I16770)
g14694(1) = NOT(I16795)
g14705(1) = NOT(I16803)
g14738(1) = NOT(I16821)
g14749(1) = NOT(I16829)
g14779(1) = NOT(I16847)
g14828(1) = NOT(I16875)
g16603(1) = NOT(I17787)
g16624(1) = NOT(I17814)
g16627(1) = NOT(I17819)
g16656(1) = NOT(I17852)
g16659(1) = NOT(I17857)
g16686(1) = NOT(I17892)
g16693(1) = NOT(I17901)
g16718(1) = NOT(I17932)
g16722(1) = NOT(I17938)
g16744(1) = NOT(I17964)
g16748(1) = NOT(I17970)
g16775(1) = NOT(I17999)
g16874(1) = NOT(I18066)
g16924(1) = NOT(I18092)
g16955(1) = NOT(I18107)
g17291(1) = NOT(I18276)
g17316(1) = NOT(I18293)
g17320(1) = NOT(I18297)
g17400(1) = NOT(I18333)
g17404(1) = NOT(I18337)
g17423(1) = NOT(I18360)
g17519(1) = NOT(I18460)
g17577(1) = NOT(I18504)
g17580(1) = NOT(I18509)
g17604(1) = NOT(I18555)
g17607(1) = NOT(I18560)
g17639(1) = NOT(I18600)
g17646(1) = NOT(I18609)
g17649(1) = NOT(I18614)
g17674(1) = NOT(I18647)
g17678(1) = NOT(I18653)
g17685(1) = NOT(I18662)
g17688(1) = NOT(I18667)
g17711(1) = NOT(I18694)
g17715(1) = NOT(I18700)
g17722(1) = NOT(I18709)
g17739(1) = NOT(I18728)
g17743(1) = NOT(I18734)
g17760(1) = NOT(I18752)
g17764(1) = NOT(I18758)
g17778(1) = NOT(I18778)
g17787(1) = NOT(I18795)
g17813(1) = NOT(I18813)
g17819(1) = NOT(I18825)
g17845(1) = NOT(I18835)
g17871(1) = NOT(I18845)
g19334(1) = NOT(I19818)
g19357(1) = NOT(I19837)
g6974(1) = NOT(I11746)
g6972(1) = NOT(I11740)
g10831(6) = NOR(g7690, g7827)
g11889(1) = NOT(g9954)
g10905(3) = NAND(g1116, g7304)
g11888(1) = NOT(g10160)
g10392(1) = NOT(g6989)
g9245(1) = NOT(I13031)
g8925(2) = NOT(I12910)
g8134(1) = NOT(I12415)
g10288(1) = NOT(I13718)
g10233(27) = NOT(I13699)
I15070(1) = NOT(g10108)
I14935(1) = NOT(g9902)
g10939(6) = NAND(g7352, g1459)
I14054(1) = NOT(g10028)
g10374(1) = NOT(g6903)
g7791(10) = NOT(I12199)
I14970(1) = NOT(g9965)
g12297(2) = NOR(g9269, g9239)
g9637(1) = NOT(I13252)
I15250(1) = NOT(g9152)
g10489(1) = NOT(g9259)
g10971(8) = NAND(g7867, g7886)
g7502(1) = NOT(I11992)
g12417(1) = NOT(g7175)
g12601(2) = NOR(g9381, g9311)
g10087(2) = NOT(I13597)
g9417(11) = NOT(I13124)
g8876(2) = NOT(I12855)
g10412(1) = NOT(g7072)
I13990(1) = NOT(g7636)
g10414(1) = NOT(g7092)
I14679(1) = NOT(g9332)
g10383(1) = NOT(g6978)
g8791(1) = NOT(I12787)
g11714(1) = NOT(g8107)
I14455(1) = NOT(g10197)
g7717(15) = NOT(I12172)
g11910(1) = NOT(g10185)
g11360(2) = NOR(g3763, g8669)
I14267(1) = NOT(g7835)
g10582(1) = NOT(g7116)
g6755(1) = NOT(I11620)
g10029(1) = NOT(I13548)
g11741(2) = NOT(g10033)
g10357(1) = NOT(g6825)
g11735(1) = NOT(g8534)
g9154(1) = NOT(I12994)
g10352(1) = NOT(g6804)
g10520(1) = NAND(g7195, g7115)
g7766(10) = NOT(I12189)
g7753(9) = NOT(I12183)
g8844(2) = NOT(I12826)
g7594(1) = NOT(I12064)
g8821(1) = NOT(I12811)
g11866(1) = NOT(g9883)
g8818(2) = NOT(I12808)
I14905(1) = NOT(g9822)
g11280(2) = NOR(g8647, g3408)
g12465(1) = NOT(g7192)
g10951(8) = NAND(g7845, g7868)
I14241(1) = NOT(g8356)
g9746(1) = NOT(I13326)
g10401(1) = NOT(g7041)
g8038(7) = NOT(I12360)
g10862(6) = NOR(g7701, g7840)
g10371(1) = NOT(g6918)
g9747(1) = NOT(I13329)
I14584(1) = NOT(g9766)
g10893(2) = NOR(g1189, g7715, g7749)
g11721(2) = NOT(g10074)
g7689(1) = NOT(I12159)
g7618(1) = NOT(I12092)
g7028(11) = NOT(I11785)
g7516(1) = NOT(I12003)
g7515(1) = NOT(I12000)
g7097(11) = NOT(I11809)
g10573(4) = NAND(g7992, g8179)
g10380(1) = NOT(g6960)
g9021(2) = NOT(I12954)
g9281(1) = NOT(I13057)
g9186(1) = NOT(I13010)
g10349(1) = NOT(g6956)
I14797(1) = NOT(g9636)
g8085(1) = NOT(I12382)
g12021(1) = NOT(g9543)
g10382(1) = NOT(g6958)
g10142(1) = NOT(I13637)
g9935(11) = NOT(I13483)
g9280(1) = NOT(I13054)
g10519(1) = NOT(g9326)
g10518(1) = NOT(g9311)
g10408(1) = NOT(g7049)
g12122(1) = NOT(g9705)
g7624(1) = NOT(I12106)
g8812(5) = NOT(I12805)
g11038(1) = NOT(g8632)
g7196(1) = NOT(I11860)
g11815(3) = NOT(g7582)
g8405(1) = NOT(I12572)
g12198(2) = NOR(g9797, g9800)
g11676(1) = NAND(g358, g8944, g376, g385)
g8032(1) = NOT(I12355)
I14033(1) = NOT(g8912)
g8974(2) = NOT(I12930)
g7994(1) = NOT(I12336)
g11884(1) = NOT(g8125)
g10399(1) = NOT(g7017)
I14967(1) = NOT(g9964)
I15223(1) = NOT(g10119)
g10415(1) = NOT(g7109)
g11110(1) = NOT(g8728)
g10664(1) = NOT(g8928)
g12729(1) = NOR(g1657, g8139)
g7566(1) = NOT(I12049)
g10356(1) = NOT(g6819)
g6867(1) = NOT(I11685)
g11607(1) = NOR(g8848, g8993, g376)
g9155(2) = NOT(I12997)
g11762(1) = NOT(g7964)
g10370(1) = NOT(g7095)
g6821(3) = NOT(I11655)
I14902(1) = NOT(g9821)
I14046(1) = NOT(g9900)
g10410(1) = NOT(g7069)
g9213(1) = NOT(I13020)
g8411(4) = NOT(I12577)
g6756(10) = NOT(I11623)
g7074(11) = NOT(I11801)
g10400(1) = NOT(g7002)
g7474(1) = NOT(I11980)
g7527(1) = NOT(I12016)
g10379(1) = NOT(g6953)
g11841(1) = NOT(g9800)
g10198(1) = NOT(I13672)
g7633(1) = NOT(I12120)
g9340(13) = NOT(I13094)
g12047(1) = NOT(g9591)
I13847(1) = NOT(g7266)
g12051(1) = NOT(g9595)
g6875(11) = NOT(I11697)
g10935(3) = NAND(g1459, g7352)
g10882(1) = NOT(g7601)
g7617(1) = NOT(I12089)
g10407(1) = NOT(g7063)
g8481(11) = NOT(I12618)
g10632(16) = AND(g7475, g7441, g890)
g10725(1) = NOT(g7846)
g7161(1) = NOT(I11843)
g7051(11) = NOT(I11793)
g10107(1) = NOT(I13606)
g12550(2) = NOR(g9300, g9259)
I14222(1) = NOT(g8286)
g10398(1) = NOT(g6999)
g10141(1) = NOT(I13634)
g10652(1) = NOT(g7601)
g9772(2) = NOT(I13352)
g9687(1) = NOT(I13287)
I15382(1) = NOT(g9071)
g10406(1) = NOT(g7046)
g10361(1) = NOT(g6841)
g8703(8) = NOT(I12709)
g12249(2) = NOR(g5763, g10096)
g8357(1) = NOT(I12538)
g10388(1) = NOT(g6983)
g7565(1) = NOT(I12046)
g10909(6) = NAND(g7304, g1116)
g11149(3) = NAND(g1564, g7948)
g10397(1) = NOT(g7018)
g7596(1) = NOT(I12070)
g10273(1) = NOT(I13708)
I14050(1) = NOT(g9963)
g12779(1) = NOT(g9444)
g12778(1) = NOT(g9856)
g7117(1) = NOT(I11816)
g10795(1) = NOT(g7202)
g12467(2) = NOR(g9472, g9407)
I15073(1) = NOT(g10109)
g10556(4) = NAND(g7971, g8133)
g12233(1) = NOT(g10338)
g11122(1) = NOT(g8751)
I14301(1) = NOT(g8571)
I15030(1) = NOT(g10073)
g10003(11) = NOT(I13539)
g11006(3) = NOR(g7686, g7836)
g6971(1) = NOT(I11737)
g11034(1) = NOT(g7611)
g10541(1) = NOT(g9407)
g6868(1) = NOT(I11688)
g10359(1) = NOT(g6830)
g10358(1) = NOT(g6827)
g12318(2) = NOR(g10172, g6451)
g7704(10) = NOT(I12167)
g10319(1) = NOT(I13740)
g11283(6) = NOR(g7953, g4991, g9064)
g11796(1) = NOT(g7985)
g8841(2) = NOT(I12823)
g8763(1) = NOT(I12749)
g10402(1) = NOT(g7023)
g6905(11) = NOT(I11708)
g7626(1) = NOT(I12112)
I14119(1) = NOT(g7824)
g8757(5) = NOT(I12746)
g11270(2) = NOR(g8431, g8434)
I14773(1) = NOT(g9581)
g8470(4) = NOT(I12605)
g10395(1) = NOT(g6995)
g11948(1) = NOT(g10224)
g12659(2) = NOR(g9451, g9392)
g6832(3) = NOT(I11665)
g6928(11) = NOT(I11716)
g8880(2) = NOT(I12861)
g8595(11) = NOT(I12666)
g10287(1) = NOT(I13715)
g8135(1) = NOT(I12418)
g7526(1) = NOT(I12013)
g7632(1) = NOT(I12117)
g10389(1) = NOT(g6986)
g8542(11) = NOT(I12644)
g10272(1) = NOT(I13705)
g12308(2) = NOR(g9951, g9954)
g6973(1) = NOT(I11743)
I15205(1) = NOT(g10139)
g9780(12) = NOT(I13360)
g8989(1) = NOT(I12935)
g10061(11) = NOT(I13581)
g7616(1) = NOT(I12086)
g7004(12) = NOT(I11777)
I14537(1) = NOT(g10106)
g7647(1) = NOT(I12132)
g10360(1) = NOT(g6836)
g10387(1) = NOT(g6996)
g8355(1) = NOT(I12534)
g11413(1) = NOT(g9100)
I14570(1) = NOT(g7932)
g12831(1) = NOT(g9569)
g9153(1) = NOT(I12991)
g10355(1) = NOT(g6816)
I14866(1) = NOT(g9748)
I14742(1) = NOT(g9534)
I13995(1) = NOT(g8744)
g10367(1) = NOT(g6870)
g10394(1) = NOT(g6994)
g8971(2) = NOT(I12927)
g7738(10) = NOT(I12176)
g10420(1) = NOT(g9239)
g9864(11) = NOT(I13424)
I14550(1) = NOT(g10072)
g11769(1) = NOT(g8626)
g10540(1) = NOT(g9392)
g10376(1) = NOT(g6923)
g10377(1) = NOT(g6940)
g8740(1) = NOT(I12735)
g12201(2) = NOR(g5417, g10047)
I14271(1) = NOT(g8456)
g11779(1) = NOT(g9602)
g10427(1) = NOT(g10053)
g10366(1) = NOT(g6895)
g10381(1) = NOT(g6957)
g11786(3) = NOT(g7549)
g10386(1) = NOT(g6982)
g10393(1) = NOT(g6991)
g10403(1) = NOT(g7040)
g8879(1) = NOT(I12858)
g11233(1) = NOT(g9664)
g11618(2) = NOR(g8114, g8070)
g9477(1) = NOT(I13149)
I14839(1) = NOT(g9689)
g11513(1) = NOT(g7948)
g10490(1) = NOT(g9274)
g9104(47) = NOT(I12987)
g12126(2) = NOR(g9989, g5069)
g10980(1) = NOT(g9051)
g11026(1) = NOT(g8434)
g12086(1) = NOT(g9654)
g11018(1) = AND(g7655, g7643, g7627)
g10354(1) = NOT(g6811)
g11326(3) = NAND(g8993, g376, g365, g370)
I15162(1) = NOT(g10176)
g10404(1) = NOT(g7026)
g12295(1) = NOT(g7139)
g12823(1) = NOT(g9206)
g11811(1) = NOT(g9724)
g8515(3) = NOT(I12631)
g10497(1) = NOT(g10102)
g11330(5) = NAND(g9483, g1193)
I13979(1) = NOT(g7733)
g7993(1) = NOT(I12333)
g11011(1) = NOT(g10274)
g12160(2) = NOR(g9721, g9724)
g10411(1) = NOT(g7086)
g12256(2) = NOR(g10136, g6105)
g10581(1) = NOT(g9529)
g7615(1) = NOT(I12083)
g12830(1) = NOT(g9995)
g10391(1) = NOT(g6988)
g10230(1) = NOT(I13694)
g10372(1) = NOT(g6900)
g9917(2) = NOT(I13473)
g11303(2) = NOR(g8497, g8500)
g6754(1) = NOT(I11617)
I14079(1) = NOT(g7231)
g8792(2) = NOT(I12790)
g7640(2) = NOT(I12128)
g7812(10) = NOT(I12214)
g11273(2) = NOR(g3061, g8620)
g6961(9) = NOT(I11734)
g11261(6) = NOR(g7928, g4801, g9030)
g6946(6) = NOT(I11721)
g7634(1) = NOT(I12123)
g10416(1) = NOT(g10318)
g11316(1) = NOT(g8967)
I14475(1) = NOT(g10175)
g12246(2) = NOR(g9880, g9883)
I14893(1) = NOT(g9819)
I14836(1) = NOT(g9688)
g11753(1) = NOT(g8587)
g11031(1) = NOT(g8609)
g11736(1) = NOT(g8165)
g11313(2) = NOR(g8669, g3759)
g10351(1) = NOT(g6802)
g6869(1) = NOT(I11691)
g12208(2) = NOR(g10096, g5759)
g9185(1) = NOT(I13007)
g10373(1) = NOT(g6917)
g11493(2) = NOR(g8964, g8967)
g11148(1) = NOR(g8052, g9197, g9174, g9050)
g11043(1) = NOT(g8561)
g11810(1) = NOT(g9664)
I14862(1) = NOT(g8092)
g6888(6) = NOT(I11701)
g12235(2) = NOR(g9234, g9206)
g8285(1) = NOT(I12497)
I14932(1) = NOT(g9901)
g10918(2) = NOR(g1532, g7751, g7778)
g8795(1) = NOT(I12793)
I14593(1) = NOT(g9978)
g10390(1) = NOT(g6987)
I14409(1) = NOT(g8364)
g11017(1) = NOT(g10289)
g11346(2) = NOR(g7980, g7964)
g10413(1) = NOT(g7110)
g8572(2) = NOT(I12654)
g8712(1) = NOT(I12712)
I14827(1) = NOT(g9686)
g11130(3) = NAND(g1221, g7918)
g10216(1) = NOT(I13684)
I14381(1) = NOT(g8300)
g11865(1) = NOT(g10124)
g12228(3) = NOR(g10222, g10206, g10184, g10335)
g8805(1) = NOT(I12799)
I14326(1) = NOT(g8607)
g11042(1) = NOT(g8691)
g12805(1) = NOT(g9511)
I14567(1) = NOT(g9708)
g11383(1) = NOT(g9061)
g11030(1) = NOT(g8292)
g6767(4) = NOT(I11626)
g12358(2) = NOR(g10019, g10022)
g11666(2) = NOR(g8172, g8125)
g6976(1) = NOT(I11750)
g7625(1) = NOT(I12109)
g7623(1) = NOT(I12103)
g10362(1) = NOT(g6850)
g8476(1) = OR(g1399, g1459, I12611)
g7593(1) = NOT(I12061)
g12082(1) = NOT(g9645)
g12345(1) = NOT(g7158)
g12399(2) = NOT(g9920)
g12804(1) = NOT(g9927)
g11415(2) = NOR(g8080, g8026)
g7595(1) = NOT(I12067)
g11563(2) = NOR(g8059, g8011)
g8922(2) = NOT(I12907)
g7542(1) = NOT(I12030)
g11306(2) = NOR(g3412, g8647)
g10409(1) = NOT(g7087)
g11012(3) = NOR(g7693, g7846)
I14999(1) = NOT(g10030)
g7148(1) = NOT(I11835)
I14505(1) = NOT(g10140)
g6772(9) = NOT(I11629)
g11385(2) = NOR(g8021, g7985)
g6856(10) = NOT(I11682)
g7121(10) = NOT(I11820)
g10621(1) = NOT(g7567)
g11252(2) = NOR(g8620, g3057)
I14896(1) = NOT(g9820)
g10564(1) = NOT(g9462)
g7586(4) = NOT(I12056)
g7660(1) = NOT(I12144)
g7659(1) = NOT(I12141)
g10872(1) = NOT(g7567)
g10405(1) = NOT(g7064)
g6977(1) = NOT(I11753)
g12440(2) = NOT(g9985)
g11214(1) = NOT(g9602)
g10350(1) = NOT(g6800)
g10396(1) = NOT(g6997)
g12170(2) = NOR(g10047, g5413)
g10378(1) = NOT(g6926)
g11991(1) = NOT(g9485)
g10881(1) = NOT(g7567)
g7648(1) = NOT(I12135)
g12708(2) = NOR(g9518, g9462)
g11849(2) = NOT(g7601)
g7674(1) = NOT(I12151)
g11374(5) = NAND(g9536, g1536)
g11833(1) = NOT(g8026)
I14158(1) = NOT(g8806)
g12738(1) = NOT(g9374)
g10897(1) = NOT(g7601)
g11812(2) = NOT(g7567)
g11033(1) = NOT(g8500)
g10369(1) = NOT(g6873)
g10368(1) = NOT(g6887)
g7543(1) = NOT(I12033)
g9478(1) = NOT(I13152)
g11344(1) = NOT(g9015)
g6782(6) = NOT(I11632)
I14823(1) = NOT(g8056)
I13968(1) = NOT(g7697)
g10808(3) = NOR(g8509, g7611)
g12088(4) = NOT(g7701)
g10615(1) = NOR(g1636, g7308)
g7558(4) = NOT(I12041)
g11927(1) = NOT(g10207)
g10428(1) = NOT(g9631)
g12361(2) = NOR(g6455, g10172)
g10375(1) = NOT(g6941)
g10323(10) = NOT(I13744)
g11357(2) = NOR(g8558, g8561)
g6789(9) = NOT(I11635)
g11832(1) = NOT(g8011)
g11861(1) = NOT(g8070)
g11083(23) = AND(g8836, g802)
g12018(1) = NOT(g9538)
g12311(2) = NOR(g6109, g10136)
g12163(2) = NOR(g5073, g9989)
g10031(1) = NOT(I13552)
g11472(1) = NOT(g7918)
g11911(1) = NOT(g10022)
g10960(1) = NOT(g9007)
g8417(1) = OR(g1056, g1116, I12583)
g11754(1) = NOT(g8229)
g10708(1) = NOT(g7836)
g7831(2) = NOT(I12227)
g12054(4) = NOT(g7690)
g8778(4) = NOT(I12758)
g6955(1) = NOT(I11726)
g12347(2) = NOR(g9321, g9274)
g12768(3) = OR(g7785, g7202)
g10353(1) = NOT(g6803)
g10295(10) = NOT(I13723)
g12752(2) = NOR(g9576, g9529)
g11171(1) = NOR(g8088, g9226, g9200, g9091)
g12419(2) = NOR(g9402, g9326)
g12015(1) = AND(g1002, g7567)
I24597(1) = AND(g5736, g5742, g9875)
g11546(1) = AND(g7289, g4375)
g11024(1) = AND(g5436, g9070)
I13937(1) = AND(g7340, g7293, g7261)
g11998(1) = NAND(g8324, g8373)
g12023(1) = NAND(g2453, g8373)
g12179(1) = AND(g9745, g10027)
g11497(1) = AND(g6398, g7192)
g11126(1) = AND(g6035, g10185)
g12186(1) = AND(g1178, g7519)
g11409(1) = NAND(g9842, g3298)
g11381(1) = NAND(g9660, g3274)
I24508(1) = AND(g9434, g9672, g5401)
g12762(4) = AND(g4358, g8977)
g10705(1) = AND(g6850, g10219, g2689)
g11834(6) = NOR(g8938, g8822)
I24600(1) = AND(g6077, g6082, g9946)
g12523(1) = NAND(g7563, g6346)
g12463(1) = NAND(g7513, g6322)
g11496(1) = AND(g4382, g7495)
g11978(2) = AND(g2629, g7462)
g11804(5) = NOR(g8938, g4975)
I24051(1) = AND(g3380, g3385, g8492)
g11019(1) = AND(g5092, g9036)
I24530(1) = AND(g9501, g9733, g5747)
g10800(1) = OR(g7517, g952)
g10822(1) = AND(g4264, g8514)
g10586(1) = NAND(g7380, g7418)
g10569(1) = NAND(g2287, g7418)
g11957(1) = NAND(g8205, g8259)
g11974(1) = NAND(g2185, g8259)
g12589(1) = NAND(g7591, g6692)
g12525(1) = NAND(g7522, g6668)
g10616(1) = AND(g7998, g174)
g10704(1) = AND(g2145, g10200, g2130)
g10999(2) = AND(g7880, g1472)
g10967(2) = AND(g7880, g1448)
g10829(1) = AND(g7289, g4375)
g11916(2) = AND(g2227, g7328)
I24075(1) = AND(g3736, g3742, g8553)
g12341(1) = NAND(g7512, g5308)
g12293(1) = NAND(g7436, g5283)
g10665(1) = AND(g209, g8292)
I13862(1) = AND(g7232, g7219, g7258)
g12521(1) = NAND(g7471, g5969)
g12356(1) = NAND(g7438, g6012)
g12307(1) = NAND(g7395, g5983)
g10796(2) = NAND(g7537, g7523)
g11491(1) = NAND(g9982, g4000)
g11445(1) = NAND(g9771, g3976)
g10568(1) = NAND(g7328, g7374)
g10552(1) = NAND(g2153, g7374)
g10675(1) = AND(g3436, g8500)
g11940(1) = NOR(g2712, g10084)
g10883(1) = AND(g3355, g9061)
g10501(1) = AND(g1233, g9007)
g11937(2) = AND(g1936, g7362)
g10726(1) = NAND(g7304, g7661, g979, g1061)
g10566(1) = NAND(g7315, g7356)
g10551(1) = NAND(g1728, g7356)
g10890(2) = AND(g7858, g1105)
g11996(1) = NAND(g7280, g2197)
g11223(1) = AND(g8281, g8505)
g11740(1) = AND(g8769, g703)
I24582(1) = AND(g9809, g9397, g6093)
g12638(1) = NAND(g7514, g6661)
g12476(1) = NAND(g7498, g6704)
g12429(1) = NAND(g7473, g6675)
g10921(1) = AND(g1548, g8685)
g12048(1) = NAND(g7369, g2040)
g10674(1) = AND(g6841, g10200, g2130)
g10732(1) = AND(g6850, g2697, g2689)
g10934(1) = AND(g9197, g7918)
I24027(1) = AND(g3029, g3034, g8426)
I24482(1) = AND(g9364, g9607, g5057)
I24552(1) = AND(g9733, g9316, g5747)
I24003(1) = AND(g8097, g8334, g3045)
g10948(2) = AND(g7880, g1478)
g10683(1) = AND(g7289, g4438)
g11116(1) = AND(g9960, g6466)
g11797(6) = NOR(g8883, g8796)
I24527(1) = AND(g9672, g9264, g5401)
I24505(1) = AND(g9607, g9229, g5057)
g11035(1) = AND(g5441, g9800)
g11142(1) = AND(g6381, g10207)
I24603(1) = AND(g9892, g9467, g6439)
g11708(1) = NAND(g10147, g10110)
g12027(1) = AND(g9499, g9729)
g10602(1) = NAND(g7411, g7451)
g10585(1) = NAND(g1996, g7451)
g10947(1) = AND(g9200, g1430)
g11950(1) = NOR(g9220, g9166)
g12346(1) = NOR(g9931, g9933)
I24549(1) = AND(g5385, g5390, g9792)
I24018(1) = AND(g8155, g8390, g3396)
g10724(1) = AND(g3689, g8728)
g10755(1) = NAND(g7352, g7675, g1322, g1404)
I24048(1) = AND(g3034, g3040, g8426)
g12466(1) = NOR(g10057, g10059)
g10898(1) = AND(g3706, g9100)
g11469(1) = NOR(g650, g9903, g645)
g10719(1) = AND(g6841, g2138, g2130)
I24625(1) = AND(g6428, g6434, g10014)
g12730(4) = AND(g9024, g4349)
g11397(1) = AND(g5360, g7139)
g11971(1) = NAND(g8249, g8302)
g11993(1) = NAND(g1894, g8302)
I24064(1) = AND(g3385, g3391, g8492)
g11047(1) = AND(g6474, g9212)
g11205(1) = AND(g8217, g8439)
g11046(1) = AND(g9889, g6120)
g12687(4) = AND(g9024, g8977)
g10902(2) = AND(g7858, g1129)
g12259(24) = AND(g9480, g640)
g11027(1) = AND(g5097, g9724)
g12043(1) = AND(g1345, g7601)
g11003(2) = AND(g7880, g1300)
g12413(1) = NAND(g7521, g5654)
g12343(1) = NAND(g7470, g5630)
g10799(1) = NOR(g347, g7541)
g11449(1) = AND(g6052, g7175)
g10925(2) = AND(g7858, g956)
I24030(1) = AND(g8390, g8016, g3396)
g11913(1) = NOR(g7197, g9166)
g12817(1) = AND(g1351, g7601)
I24054(1) = AND(g8443, g8075, g3747)
I24015(1) = AND(g8334, g7975, g3045)
g10625(1) = AND(g3431, g7926)
g10699(4) = NOR(g8526, g1514)
g10610(1) = NAND(g7462, g7490)
g10605(1) = NAND(g2555, g7490)
I24524(1) = AND(g5041, g5046, g9716)
g11443(1) = NAND(g9916, g3649)
g11411(1) = NAND(g9713, g3625)
g10803(1) = NOR(g1384, g7503)
g12591(1) = NOR(g504, g9040)
I24616(1) = AND(g6082, g6088, g9946)
g12587(1) = NAND(g7497, g6315)
g12428(1) = NAND(g7472, g6358)
g12357(1) = NAND(g7439, g6329)
g10707(1) = AND(g3787, g8561)
g12411(1) = NAND(g7393, g5276)
g12244(1) = NAND(g7343, g5320)
g12197(1) = NAND(g7296, g5290)
g12065(1) = AND(g9557, g9805)
g12234(1) = NOR(g9776, g9778)
I24555(1) = AND(g9559, g9809, g6093)
g10793(1) = NOR(g1389, g7503)
g10917(1) = AND(g9174, g1087)
g12219(1) = AND(g1189, g7532)
g10706(1) = AND(g3338, g8691)
g10624(1) = AND(g8387, g3072)
g10709(1) = NOR(g7499, g351)
g11891(1) = NOR(g812, g9166)
g10802(1) = OR(g7533, g1296)
g11960(2) = AND(g2495, g7424)
g10655(1) = AND(g8440, g3423)
g11244(1) = AND(g8346, g8566)
I24585(1) = AND(g9621, g9892, g6439)
I24576(1) = AND(g5390, g5396, g9792)
g10619(1) = AND(g3080, g7907)
g11967(1) = AND(g311, g7802)
g11010(1) = AND(g4698, g8933)
g10677(1) = AND(g4141, g7611)
I14198(1) = AND(g225, g8237, g232, g8180)
g10676(1) = AND(g8506, g3774)
g11201(1) = NOR(g4125, g7765)
g10654(1) = AND(g3085, g8434)
g11023(1) = AND(g9669, g5084)
g10878(2) = AND(g7858, g1135)
g12284(1) = AND(g1532, g7557)
I24067(1) = AND(g3731, g3736, g8553)
g10584(1) = NAND(g7362, g7405)
g10567(1) = NAND(g1862, g7405)
g11016(1) = AND(g4888, g8984)
g12019(1) = NAND(g7322, g1906)
g11893(2) = AND(g1668, g7268)
g11543(1) = NAND(g9714, g3969)
g11424(1) = NAND(g9662, g4012)
g11395(1) = NAND(g9601, g3983)
g10666(4) = NOR(g8462, g1171)
g10841(9) = AND(g8509, g8567)
g11939(2) = AND(g2361, g7380)
g11953(1) = NAND(g8195, g8241)
g11970(1) = NAND(g1760, g8241)
g12761(1) = AND(g969, g7567)
g10604(1) = NAND(g7424, g7456)
g10587(1) = NAND(g2421, g7456)
g10720(1) = AND(g2704, g10219, g2689)
g12052(1) = NAND(g7387, g2465)
I24033(1) = AND(g8219, g8443, g3747)
g10684(1) = AND(g7998, g411)
g11915(2) = AND(g1802, g7315)
g11037(1) = AND(g6128, g9184)
I24546(1) = AND(g5046, g5052, g9716)
g10760(1) = NOR(g1046, g7479)
g10873(1) = AND(g3004, g9015)
g11036(1) = AND(g9806, g5774)
g12135(1) = AND(g9684, g9959)
g11975(1) = NAND(g8267, g8316)
g11997(1) = NAND(g2319, g8316)
I14225(1) = AND(g8457, g255, g8406, g262)
g10565(1) = AND(g8182, g424)
g11934(1) = NAND(g8139, g8187)
g11952(1) = NAND(g1624, g8187)
g11994(1) = NAND(g8310, g8365)
g12020(1) = NAND(g2028, g8365)
g12812(4) = AND(g518, g9158)
g12795(1) = AND(g1312, g7601)
g11370(1) = OR(g8807, g550)
g10550(1) = NAND(g7268, g7308)
g10529(1) = NAND(g1592, g7308)
I24579(1) = AND(g5731, g5736, g9875)
g11780(5) = NOR(g4899, g8822)
g11969(1) = NAND(g7252, g1636)
g11755(5) = NOR(g4709, g8796)
g10820(1) = NAND(g9985, g9920, g9843)
g11115(1) = AND(g6133, g9954)
g12296(1) = NOR(g9860, g9862)
g12794(1) = AND(g1008, g7567)
g11489(1) = NAND(g9661, g3618)
g11394(1) = NAND(g9600, g3661)
g11356(1) = NAND(g9552, g3632)
g12418(1) = NOR(g9999, g10001)
g12099(1) = AND(g9619, g9888)
g11384(1) = NOR(g8538, g8540)
g11441(1) = NAND(g9599, g3267)
g11355(1) = NAND(g9551, g3310)
g11302(1) = NAND(g9496, g3281)
g10827(1) = AND(g8914, g4258)
g12220(1) = AND(g1521, g7535)
g11114(1) = AND(g5689, g10160)
g11773(5) = NOR(g8883, g4785)
g11414(1) = NOR(g8591, g8593)
I24619(1) = AND(g6423, g6428, g10014)
g10998(1) = AND(g8567, g8509, g8451, g7650)
g11992(1) = NAND(g7275, g1772)
g11345(1) = NOR(g8477, g8479)
g11163(1) = AND(g6727, g10224)
g10896(1) = AND(g1205, g8654)
g11932(1) = NOR(g843, g9166)
g11029(1) = AND(g5782, g9103)
g11028(1) = AND(g9730, g5428)
g12527(10) = AND(g8680, g667)
g10626(1) = AND(g4057, g7927)
g12022(1) = NAND(g7335, g2331)
g10856(1) = AND(g4269, g8967)
g11045(1) = AND(g5787, g9883)
g10736(1) = AND(g4040, g8751)
g10528(1) = AND(g1576, g9051)
g12459(1) = NAND(g7437, g5623)
g12306(1) = NAND(g7394, g5666)
g12245(1) = NAND(g7344, g5637)
g12369(1) = NAND(g9049, g637)
g10657(1) = AND(g8451, g4064)
g10801(1) = NOR(g1041, g7479)
g10970(1) = AND(g854, g9582)
g11044(1) = AND(g5343, g10124)
g12087(1) = NAND(g7431, g2599)
g11427(1) = AND(g5706, g7158)
g11366(1) = AND(g5016, g10338)
g12461(1) = NAND(g7536, g6000)
g12415(1) = NAND(g7496, g5976)
g10656(1) = AND(g3782, g7952)
g12024(1) = NAND(g8381, g8418)
g12053(1) = NAND(g2587, g8418)
g11127(1) = AND(g6479, g10022)
g10966(1) = AND(g9226, g7948)
g11956(2) = AND(g2070, g7411)
g11999(1) = NOR(g9654, g7423)
g12025(1) = NOR(g9705, g7461)
g8921(1) = OR(I12902, I12903)
g10821(1) = NOR(g7503, g1384)
g8790(1) = OR(I12782, I12783)
g10511(3) = NAND(g4628, g7202, g4621)
g11184(1) = NOR(g513, g9040)
g11958(1) = NOR(g9543, g7327)
g11380(1) = OR(g8583, g8530)
g11976(1) = NOR(g9595, g7379)
g11995(1) = NOR(g9645, g7410)
g11972(1) = NOR(g9591, g7361)
g11213(1) = NOR(g4776, g7892, g9030)
g11191(1) = NOR(g4776, g4801, g9030)
g11935(1) = NOR(g9485, g7267)
g11232(1) = NOR(g4966, g7898, g9064)
g11203(1) = NOR(g4966, g4991, g9064)
g11954(1) = NOR(g9538, g7314)
g10819(1) = NOR(g7479, g1041)
g11566(4) = NOR(g3161, g7964)
g11435(5) = NOR(g8107, g3171)
g12169(1) = NAND(g9804, g5448)
I13443(1) = NAND(g262, I13442)
I14185(2) = NAND(g8442, g3470)
I14516(2) = NAND(g10147, g661)
I12346(1) = NAND(g3111, I12344)
I14883(2) = NAND(g9500, g5489)
g11426(1) = NAND(g8742, g4878)
g11190(1) = NAND(g8539, g3447)
I15087(2) = NAND(g9832, g2393)
g12084(1) = NAND(g2342, g8211)
I13391(1) = NAND(g1821, I13390)
I13392(1) = NAND(g1825, I13390)
I11865(1) = NAND(g4434, I11864)
I11866(1) = NAND(g4401, I11864)
I13510(1) = NAND(g2089, I13509)
I13511(1) = NAND(g2093, I13509)
g12323(8) = NAND(g9480, g640)
g11968(1) = NAND(g837, g9334, g9086)
g10922(2) = NOR(g7650, g4057)
I13110(1) = NAND(g5808, I13109)
g12000(1) = NAND(g8418, g2610)
g11312(1) = NAND(g8565, g3794)
g10715(3) = NOR(g8526, g8466)
g11707(1) = NAND(g8718, g4864)
I14609(2) = NAND(g8993, g8678)
g11979(1) = NAND(g9861, g5452)
g12639(1) = NAND(g10194, g6682, g6732)
I12288(1) = NAND(g1484, I12287)
I12289(1) = NAND(g1300, I12287)
g11747(5) = NOR(g3530, g8114)
g12416(1) = NAND(g10133, g7064, g10166)
g10617(1) = NAND(g10151, g9909)
I12252(1) = NAND(g1124, I12251)
g12553(4) = NOR(g5170, g9206)
g12014(1) = NAND(g7197, g703)
g11658(4) = NOR(g8021, g3506)
g11527(5) = NOR(g8165, g8114)
g10623(1) = NAND(g10181, g9976)
I13751(1) = NAND(g4584, I13749)
g12755(4) = NOR(g6555, g9407)
g10491(5) = NOR(g6573, g9576)
g12116(1) = NAND(g2051, g8255)
g12680(5) = NOR(g9631, g9576)
g12632(5) = NOR(g9631, g6565)
g11715(4) = NOR(g8080, g8026)
g11537(5) = NOR(g8229, g3873)
g11846(2) = NOR(g7635, g7518, g7548)
g12340(1) = NAND(g4888, g8984)
g12035(1) = NAND(g10000, g6144)
g11692(4) = NOR(g8021, g7985)
I15298(2) = NAND(g10112, g1982)
I13402(1) = NAND(g2246, I13401)
I13403(1) = NAND(g2250, I13401)
I12205(1) = NAND(g1135, I12203)
g10759(1) = NAND(g7537, g324)
g11679(6) = NAND(g8836, g802)
g10421(5) = NOR(g6227, g9518)
I14991(2) = NAND(g9685, g6527)
g11933(1) = NAND(g837, g9334, g7197)
g11951(1) = NAND(g9166, g847, g703)
g12222(1) = NAND(g8310, g2028)
g11653(4) = NOR(g7980, g7964)
g11729(5) = NOR(g3179, g8059)
g12117(2) = NOR(g10113, g9755)
I14204(2) = NAND(g8508, g3821)
I15306(2) = NAND(g10116, g2407)
g10695(3) = NOR(g8462, g8407)
I15340(2) = NAND(g10154, g2541)
g12604(4) = NOR(g5517, g9239)
g12798(5) = NOR(g5535, g9381)
g11610(4) = NOR(g7980, g3155)
I13044(1) = NAND(g5115, I13043)
I13045(1) = NAND(g5120, I13043)
g12700(4) = NOR(g9321, g5857)
g12515(5) = NOR(g9511, g5873)
I15333(2) = NAND(g10152, g2116)
I13519(1) = NAND(g2514, I13518)
I13520(1) = NAND(g2518, I13518)
g11119(2) = NOR(g9180, g9203)
g11279(1) = NAND(g8504, g3443)
g12317(1) = NAND(g10026, g6486)
g12073(1) = NAND(g10058, g6490)
g11669(4) = NOR(g3863, g8026)
g12374(2) = NOR(g2185, g8205)
g12255(1) = NAND(g9958, g6140)
I11825(1) = NAND(g4593, I11824)
I11826(1) = NAND(g4601, I11824)
g12464(1) = NAND(g10169, g7087, g10191)
g12797(1) = NAND(g10275, g7655, g7643, g7627)
g12113(2) = NOR(g1648, g8187)
I12204(1) = NAND(g1094, I12203)
g12292(1) = NAND(g4698, g8933)
I13140(1) = NAND(g6154, I13139)
I13141(1) = NAND(g6159, I13139)
g12153(1) = NAND(g2610, g8330)
g12193(2) = NOR(g2342, g8316)
g12780(4) = NOR(g9402, g9326)
I13444(1) = NAND(g239, I13442)
I13453(1) = NAND(g1955, I13452)
g12154(2) = NOR(g10155, g9835)
I13111(1) = NAND(g5813, I13109)
I15363(2) = NAND(g10182, g2675)
I12402(1) = NAND(g3808, I12401)
I12403(1) = NAND(g3813, I12401)
g12526(1) = NAND(g10194, g7110, g10213)
I12373(1) = NAND(g3457, I12372)
I12374(1) = NAND(g3462, I12372)
g10622(1) = NAND(g10178, g9973)
g12460(1) = NAND(g10093, g5644, g5694)
g12344(1) = NAND(g10093, g7041, g10130)
I13565(1) = NAND(g2648, I13564)
I13464(1) = NAND(g2384, I13462)
g10653(1) = NAND(g10204, g10042)
g11584(5) = NOR(g8229, g8172)
I14788(2) = NAND(g9891, g6167)
g12042(1) = NAND(g9086, g703)
g11990(1) = NAND(g9166, g703)
g11892(1) = NAND(g7777, g9086)
g12150(2) = NOR(g2208, g8259)
I14289(2) = NAND(g8282, g3835)
g11936(1) = NAND(g8241, g1783)
g12192(1) = NAND(g8267, g2319)
g10609(1) = NAND(g10111, g9826)
I12097(1) = NAND(g1339, I12096)
g12522(1) = NAND(g10133, g5990, g6040)
I13750(1) = NAND(g4608, I13749)
g12824(5) = NOR(g5881, g9451)
I12850(1) = NAND(g4277, I12848)
g11396(1) = NAND(g8713, g4688)
g11674(1) = NAND(g8676, g4674)
g11117(1) = NAND(g8087, g8186, g8239)
g10598(2) = NAND(g7191, g6404)
g12739(4) = NOR(g9321, g9274)
g12662(4) = NOR(g5863, g9274)
I15121(2) = NAND(g9910, g2102)
g12651(4) = NOR(g9269, g5511)
g10899(2) = NOR(g4064, g8451)
g11639(1) = NAND(g8933, g4722)
I13383(1) = NAND(g269, I13382)
I13384(1) = NAND(g246, I13382)
g10515(2) = NAND(g10337, g5022)
I12730(1) = NAND(g4287, I12728)
I12241(1) = NAND(g1111, I12240)
I12242(1) = NAND(g1105, I12240)
g12050(2) = NOR(g10038, g9649)
I12877(1) = NAND(g4200, I12876)
I12878(1) = NAND(g4180, I12876)
g11442(1) = NAND(g8644, g3288, g3343)
I13183(1) = NAND(g6500, I13182)
g12443(5) = NOR(g9374, g9300)
g12483(2) = NOR(g2453, g8324)
I14247(2) = NAND(g1322, g8091)
I15041(2) = NAND(g9752, g1834)
I13850(2) = NAND(g862, g7397)
g12453(5) = NOR(g9444, g5527)
g12008(1) = NAND(g9932, g5798)
g12152(1) = NAND(g2485, g8324)
g12081(2) = NOR(g10079, g9694)
I14764(2) = NAND(g9808, g5821)
I15128(2) = NAND(g9914, g2527)
g12085(2) = NOR(g10082, g9700)
g12405(5) = NOR(g9374, g5180)
g11697(4) = NOR(g8080, g3857)
g12744(4) = NOR(g9402, g6203)
g12581(5) = NOR(g9569, g6219)
I13731(1) = NAND(g4537, I13729)
I15253(2) = NAND(g10078, g1848)
g11039(2) = NOR(g9056, g9092)
I15174(2) = NAND(g9977, g2661)
g11251(1) = NAND(g8438, g3092)
g11483(5) = NOR(g8165, g3522)
I15262(2) = NAND(g10081, g2273)
I12271(1) = NAND(g956, I12269)
g11869(2) = NOR(g7649, g7534, g7581)
g11490(1) = NAND(g8666, g3639, g3694)
g11412(1) = NAND(g8666, g6918, g8697)
g12785(4) = NOR(g9472, g6549)
g11881(2) = NAND(g9060, g3361)
g12432(2) = NOR(g1894, g8249)
g11320(2) = NAND(g4633, g4621, g7202)
I14955(2) = NAND(g9620, g6181)
g11945(2) = NOR(g7212, g7228)
g10946(1) = NAND(g1489, g7876)
I13335(1) = NAND(g1687, I13334)
I13336(1) = NAND(g1691, I13334)
g11885(2) = NOR(g7153, g7167)
g12149(1) = NAND(g8205, g2185)
I14480(2) = NAND(g10074, g655)
g12148(1) = NAND(g2060, g8310)
I12545(1) = NAND(g191, I12544)
I13184(1) = NAND(g6505, I13182)
g12412(1) = NAND(g10044, g5297, g5348)
g12695(4) = NOR(g9269, g9239)
I12546(1) = NAND(g194, I12544)
g12593(4) = NOR(g9234, g5164)
g12772(5) = NOR(g5188, g9300)
g12112(1) = NAND(g8139, g1624)
g12333(2) = NOR(g1624, g8139)
I13454(1) = NAND(g1959, I13452)
I14853(2) = NAND(g9433, g5142)
g12017(2) = NOR(g9969, g9586)
I15212(2) = NAND(g10035, g1714)
I12842(1) = NAND(g4235, I12840)
I14712(2) = NAND(g9671, g5128)
I13730(1) = NAND(g4534, I13729)
I14257(2) = NAND(g8154, g3133)
I15051(2) = NAND(g9759, g2259)
I14816(2) = NAND(g9962, g6513)
g12232(1) = NAND(g8804, g4878)
g12223(2) = NOR(g2051, g8365)
g12288(2) = NOR(g2610, g8418)
g10649(2) = NOR(g1183, g8407)
I12270(1) = NAND(g1141, I12269)
I14733(2) = NAND(g9732, g5475)
g12622(5) = NOR(g9569, g9518)
g11763(5) = NOR(g3881, g8172)
I12219(1) = NAND(g1478, I12217)
g12806(4) = NOR(g9472, g9407)
g11020(2) = NAND(g9187, g9040)
g12080(1) = NAND(g1917, g8201)
I12218(1) = NAND(g1437, I12217)
g12226(2) = NOR(g2476, g8373)
I14923(2) = NAND(g9558, g5835)
g12145(1) = NAND(g8195, g1760)
g10671(2) = NOR(g1526, g8466)
I12470(1) = NAND(g392, I12468)
g10884(2) = NOR(g7650, g8451)
I13499(1) = NAND(g232, I13497)
g12711(4) = NOR(g6209, g9326)
I12075(1) = NAND(g996, I12074)
I13498(1) = NAND(g255, I13497)
g12225(1) = NAND(g8324, g2453)
I15002(2) = NAND(g9691, g1700)
g12571(5) = NOR(g9511, g9451)
g11961(1) = NAND(g9777, g5105)
g12079(1) = NAND(g1792, g8195)
g12078(1) = NAND(g8187, g8093)
I11879(1) = NAND(g4430, I11877)
g11675(1) = NAND(g8984, g4912)
I11878(1) = NAND(g4388, I11877)
g12159(1) = NAND(g8765, g4864)
g12125(1) = NAND(g9728, g5101)
g10583(1) = NAND(g7475, g862)
I13079(1) = NAND(g5467, I13077)
I13078(1) = NAND(g5462, I13077)
I14169(2) = NAND(g8389, g3119)
g12289(2) = NAND(g9978, g9766, g9708)
g12646(4) = NOR(g9234, g9206)
g11959(1) = NAND(g8316, g2342)
g11172(1) = NAND(g8478, g3096)
I12729(1) = NAND(g4291, I12728)
I12098(1) = NAND(g1322, I12096)
I12345(1) = NAND(g3106, I12344)
g12195(1) = NAND(g2619, g8381)
g12540(2) = NOR(g2587, g8381)
g12016(1) = NAND(g1648, g8093)
g12121(2) = NOR(g10117, g9762)
g12437(2) = NOR(g2319, g8267)
g11002(1) = NAND(g7475, g862)
g12188(1) = NAND(g8249, g1894)
g12124(1) = NAND(g8741, g4674)
g11245(2) = NAND(g7636, g7733, g7697)
g12294(1) = NAND(g10044, g7018, g10090)
I14228(2) = NAND(g979, g8055)
I14508(2) = NAND(g370, g8721)
g11382(1) = NAND(g8644, g6895, g8663)
g11473(5) = NOR(g8107, g8059)
I15078(2) = NAND(g9827, g1968)
g12505(5) = NOR(g9444, g9381)
I14275(2) = NAND(g8218, g3484)
g12822(1) = NAND(g6978, g7236, g7224, g7163)
g10916(1) = NAND(g1146, g7854)
g12194(1) = NAND(g8373, g8273)
g11544(1) = NAND(g8700, g3990, g4045)
g11446(1) = NAND(g8700, g6941, g8734)
g12588(1) = NAND(g10169, g6336, g6386)
I12469(1) = NAND(g405, I12468)
g12196(1) = NAND(g8764, g4688)
g12119(1) = NAND(g2351, g8267)
g12118(1) = NAND(g8259, g8150)
g11200(1) = NAND(g8592, g3798)
g11955(1) = NAND(g8302, g1917)
g11621(4) = NOR(g3512, g7985)
g10618(1) = NAND(g10153, g9913)
I14350(2) = NAND(g8890, g8848)
g12111(1) = NAND(g847, g9166)
I12278(1) = NAND(g1467, I12277)
I12279(1) = NAND(g1472, I12277)
I12849(1) = NAND(g4281, I12848)
g10601(1) = NAND(g896, g7397)
I12841(1) = NAND(g4222, I12840)
I12263(1) = NAND(g1448, I12261)
g10537(2) = NAND(g7138, g5366)
g12185(1) = NAND(g9905, g799)
g11977(1) = NAND(g8373, g2476)
g11858(2) = NAND(g9014, g3010)
g12083(1) = NAND(g2217, g8205)
g12046(2) = NOR(g10036, g9640)
I13566(1) = NAND(g2652, I13564)
g10928(1) = NAND(g8181, g8137, g417)
g12115(1) = NAND(g1926, g8249)
g10578(2) = NAND(g7174, g6058)
g11938(1) = NAND(g8259, g2208)
g12371(2) = NOR(g1760, g8195)
g12207(1) = NAND(g9887, g5794)
I12262(1) = NAND(g1454, I12261)
g11155(4) = NAND(g4776, g7892, g9030)
g12114(1) = NAND(g8241, g8146)
g10614(1) = NAND(g9024, g8977, g8928)
g12049(1) = NAND(g2208, g8150)
g11914(1) = NAND(g8187, g1648)
g10561(2) = NAND(g7157, g5712)
g11924(2) = NOR(g7187, g7209)
I13463(1) = NAND(g2380, I13462)
I12076(1) = NAND(g979, I12074)
g11973(1) = NAND(g8365, g2051)
g12045(1) = NAND(g1783, g8146)
g10929(4) = NAND(g1099, g7854)
g12147(1) = NAND(g8302, g8201)
g12151(1) = NAND(g8316, g8211)
g12227(1) = NAND(g8418, g8330)
g12044(1) = NAND(g1657, g8139)
g12120(1) = NAND(g2476, g8273)
g10961(4) = NAND(g1442, g7876)
g11216(1) = NOR(g7998, g8037)
g12189(2) = NOR(g1917, g8302)
g12146(2) = NOR(g1783, g8241)
g11173(4) = NAND(g4966, g7898, g9064)
g12190(1) = NAND(g8365, g8255)
g11231(1) = NOR(g7928, g4801, g4793)
g11907(2) = NOR(g7170, g7184)
g11134(1) = NAND(g8138, g8240, g8301)
g10603(1) = NAND(g10077, g9751)
g11903(2) = NAND(g9099, g3712)
g11862(2) = NOR(g7134, g7150)
I13066(1) = NAND(g4308, I13065)
I13067(1) = NAND(g4304, I13065)
g12479(2) = NOR(g2028, g8310)
g10611(1) = NAND(g10115, g9831)
g11107(2) = NOR(g9095, g9177)
g11248(1) = NOR(g7953, g4991, g4983)
g12287(1) = NAND(g8381, g2587)
I12253(1) = NAND(g1129, I12251)
g12486(1) = NOR(g9055, g9013, g8957, g8905)
g12252(2) = NOR(g9995, g10185)
g12166(2) = NOR(g9856, g10124)
g12821(1) = NOR(g7132, g10223, g7149, g10261)
g10555(1) = NOR(g7227, g4601, g4608)
g11363(2) = NOR(g8626, g8751)
g12204(2) = NOR(g9927, g10160)
g12364(2) = NOR(g10102, g10224)
g10510(1) = NOR(g7183, g4593, g4584)
g11309(2) = NOR(g8587, g8728)
g12314(2) = NOR(g10053, g10207)
g12435(1) = NOR(g9012, g8956, g8904, g8863)
g11276(2) = NOR(g8534, g8691)
g13297(1) = NOT(g10831)
g13103(1) = NOT(g10905)
g12884(1) = NOT(g10392)
g11181(1) = NOT(g8134)
g10571(1) = NOT(g10233)
g14339(2) = NOR(g12289, g2735)
g12217(1) = NOT(I15070)
I14749(1) = NOT(g10031)
g13190(1) = NOT(g10939)
g10816(2) = NOT(I14054)
g13134(2) = NAND(g11134, g8470)
g12110(1) = NOT(I14970)
g12922(1) = NOT(g12297)
g12321(1) = NOT(g9637)
g14981(2) = NAND(g12785, g12632)
g14782(2) = NAND(g12755, g10491)
g14933(2) = NAND(g12700, g12571)
g12381(17) = NOT(I15223)
g12450(2) = NAND(g7738, g10281)
I14833(1) = NOT(g10142)
g13625(1) = NOT(g10971)
g14848(2) = NAND(g12651, g12453)
g11250(1) = NOT(g7502)
g12936(1) = NOT(g12601)
I16231(1) = NOT(g10520)
g10830(1) = NOT(g10087)
I14653(1) = NOT(g9417)
I14671(1) = NOT(g7717)
g13990(2) = NAND(g11669, g11584)
g10430(41) = NOT(I13847)
g14098(2) = NAND(g11566, g8864)
g12909(1) = NOT(g10412)
g12543(2) = NOT(g9417)
g14691(2) = NAND(g12695, g12505)
g10678(4) = NOT(I13990)
g12908(1) = NOT(g10414)
g11867(1) = NOT(I14679)
I14702(1) = NOT(g7717)
I14576(1) = NOT(g8791)
g11450(16) = NOT(I14455)
g11819(1) = NOT(g7717)
g11048(34) = NOT(I14158)
g13707(1) = NOT(g11360)
g11202(1) = NOT(I14267)
I16917(1) = NOT(g10582)
g11988(1) = NOT(I14836)
I13762(1) = NOT(g6755)
g11984(1) = NOT(g9186)
I14830(1) = NOT(g10141)
g14665(2) = NAND(g12604, g12798)
I14745(1) = NOT(g10029)
g12841(1) = NOT(g10357)
g10981(16) = NOT(I14119)
g12835(1) = NOT(g10352)
I14761(1) = NOT(g7753)
g14011(2) = NAND(g10295, g11473)
g11402(1) = NOT(g7594)
g14918(2) = NAND(g12646, g12772)
g12933(2) = NAND(g7150, g10515)
g10419(1) = NOT(g8821)
I14727(1) = NOT(g7753)
g10418(1) = NOT(g8818)
g12041(1) = NOT(I14905)
g12430(1) = NOT(I15250)
I14579(1) = NOT(g8792)
g13706(1) = NOT(g11280)
g13756(4) = NAND(g203, g12812)
g13260(3) = NAND(g1116, g10666)
g13624(1) = NOT(g10951)
g12640(1) = NOT(I15382)
g11432(2) = NAND(g10295, g8864)
g13885(1) = NOT(g10862)
g13763(1) = NOT(g10971)
g13284(2) = NAND(g10695, g1157)
g12863(1) = NOT(g10371)
g14943(2) = NAND(g7791, g12622)
g14797(2) = NAND(g12593, g12405)
g13314(1) = NOT(g10893)
g13596(1) = NOT(g10971)
g11431(1) = NOT(g7618)
g12402(2) = NAND(g7704, g10266)
g14953(2) = NAND(g12646, g12405)
g14974(2) = NAND(g12744, g12622)
g11269(1) = NOT(g7516)
g12760(1) = NOT(g10272)
g11268(1) = NOT(g7515)
g12790(2) = NOT(g7097)
g14817(2) = NAND(g12711, g12622)
g13655(1) = NOT(g10573)
g12873(1) = NOT(g10380)
g10570(1) = NOT(g9021)
g11930(1) = NOT(g9281)
g12143(1) = NOT(I14999)
g12834(1) = NOT(g10349)
g11965(1) = NOT(I14797)
g10823(3) = AND(g7704, g5180, g5188)
g12614(7) = NOT(g9935)
g14157(2) = NAND(g11715, g11763)
g12905(1) = NOT(g10408)
g10738(2) = NAND(g6961, g10308)
g11204(1) = NOT(I14271)
g11468(1) = NOT(g7624)
g13861(3) = NAND(g1459, g10671)
g11677(1) = NOT(g7689)
g14048(2) = NAND(g11658, g11483)
g14215(1) = NOT(g12198)
I15937(1) = NOT(g11676)
g11143(1) = NOT(g8032)
g10588(1) = AND(g7004, g5297)
g10887(2) = AND(g7812, g6565, g6573)
g12891(1) = NOT(g10399)
g11928(1) = NOT(I14742)
g12109(1) = NOT(I14967)
I14964(1) = NOT(g10230)
g14627(2) = NAND(g12553, g12772)
I15800(1) = NOT(g11607)
g14773(2) = NAND(g12711, g12581)
I16747(1) = NOT(g12729)
g11373(1) = NOT(g7566)
g12840(1) = NOT(g10356)
g14864(2) = NAND(g7791, g10421)
g13898(2) = NAND(g11621, g11747)
g14861(2) = NAND(g12744, g10341)
g10554(1) = NOT(g8974)
g10608(1) = NOT(g9155)
g11964(1) = NOT(g9154)
g11985(1) = NOT(I14827)
g13216(1) = NOT(g10939)
g12862(1) = NOT(g10370)
g15033(2) = NAND(g12806, g7142)
g13923(2) = NAND(g11692, g11527)
g13330(2) = NAND(g4664, g11006)
g12040(1) = NOT(I14902)
g10805(2) = NOT(I14046)
g12904(1) = NOT(g10410)
g13569(1) = NOT(g10951)
g10761(1) = NOT(g8411)
g11129(1) = NOT(g7994)
I15033(1) = NOT(g10273)
I14623(1) = NOT(g8925)
g14130(2) = NAND(g11621, g8906)
g11293(1) = NOT(g7527)
g12872(1) = NOT(g10379)
I14899(1) = NOT(g10198)
g11510(1) = NOT(g7633)
I14633(1) = NOT(g9340)
g11615(2) = NOT(g6875)
g13116(1) = NOT(g10935)
g14021(2) = NAND(g11697, g8958)
I14589(1) = NOT(g8818)
g14151(2) = NAND(g11692, g11483)
I13872(1) = NOT(g7474)
g11430(1) = NOT(g7617)
g12820(1) = NOT(g10233)
I14305(1) = NOT(g8805)
g14841(2) = NAND(g12593, g12443)
g13142(1) = NOT(g10632)
g12929(1) = NOT(g12550)
g11165(1) = NOT(I14222)
g12578(2) = NAND(g7791, g10341)
g13202(6) = NOR(g8347, g10511)
g10804(1) = NOT(g9772)
g10590(6) = AND(g7246, g7392, I13937)
g14406(1) = NOT(g12249)
g11236(1) = NOT(g8357)
g11405(3) = NAND(g2741, g2735, g6856, g2748)
g12881(1) = NOT(g10388)
g13175(1) = NOT(g10909)
g10498(1) = NOT(g7161)
I14630(1) = NOT(g7717)
g14004(1) = NOT(g11149)
g15024(2) = NAND(g12780, g10421)
g10613(1) = NOT(g10233)
g12890(1) = NOT(g10397)
g11164(1) = NOT(g8085)
g13209(1) = NOT(g10632)
g10812(2) = NOT(I14050)
g13980(2) = NAND(g10295, g11435)
g12945(1) = NOT(g12467)
g14776(2) = NAND(g12780, g12622)
g14727(2) = NAND(g12604, g12505)
g14895(2) = NAND(g7766, g12571)
g11989(1) = NOT(I14839)
g12641(2) = AND(g10295, g3171, g3179)
g13593(1) = NOT(g10556)
g12182(1) = NOT(I15030)
g12672(7) = NOT(g10003)
g13565(1) = NOT(g11006)
g12911(2) = OR(g10278, g12768)
g14915(2) = NAND(g12553, g10266)
g15014(2) = NAND(g12785, g12680)
I13857(1) = NOT(g9780)
g12897(1) = NOT(g10400)
g14908(2) = NAND(g7812, g10491)
I13779(1) = NOT(g6868)
I14192(1) = NOT(g10233)
g14535(1) = NOT(g12318)
g13342(2) = NOR(g10961, g10935)
g10364(1) = NOT(g6869)
g14058(2) = NAND(g7121, g11537)
g12076(1) = NOT(g9280)
g12811(1) = NOT(g10319)
g14029(1) = NOT(g11283)
g14656(2) = NAND(g12553, g12405)
g14008(2) = NAND(g11610, g11435)
g10741(12) = NOT(g8411)
g10429(1) = NOT(g7148)
g12896(1) = NOT(g10402)
g14905(2) = NAND(g12785, g7142)
g14984(2) = NAND(g7812, g12680)
g13307(3) = NAND(g1116, g10695)
g11192(1) = NOT(g8038)
g11663(2) = NOT(g6905)
g13663(1) = NOT(g10971)
g14234(2) = NAND(g9177, g11881)
g14258(2) = NAND(g9203, g11903)
g13483(1) = NOT(g11270)
g11215(1) = NOT(g8285)
g12378(2) = NOT(g9417)
g11949(1) = NOT(I14773)
g10794(1) = NOT(g8470)
g14223(2) = NAND(g9092, g11858)
g10838(2) = AND(g7738, g5527, g5535)
g12944(1) = NOT(g12659)
g11702(2) = NOT(g6928)
g11182(1) = NOT(I14241)
g13621(1) = NOT(g10573)
g12793(1) = NOT(g10287)
I14644(1) = NOT(g7717)
g11183(1) = NOT(g8135)
g14041(2) = NAND(g11610, g11473)
g11509(1) = NOT(g7632)
g10612(1) = NOT(g10233)
I14684(1) = NOT(g7717)
g13121(2) = NAND(g11117, g8411)
g14813(2) = NAND(g7766, g12824)
g15018(2) = NAND(g12739, g12515)
g14251(1) = NOT(g12308)
I13802(1) = NOT(g6971)
I16024(1) = NOT(g11171)
g11912(1) = NOT(g8989)
g11592(14) = NOT(I14537)
g12880(1) = NOT(g10387)
g11691(1) = NOT(I14570)
g10776(16) = NOT(I14033)
g12629(2) = NAND(g7812, g7142)
g13960(2) = NAND(g11669, g11537)
g12887(1) = NOT(g10394)
g11640(11) = NOT(I14550)
g12843(1) = NOT(g10359)
g14879(2) = NAND(g12646, g10266)
g12869(1) = NOT(g10376)
g14914(1) = NOR(g12822, g12797)
g12868(1) = NOT(g10377)
g10542(1) = NOT(g7196)
g14377(1) = NOT(g12201)
I14660(1) = NOT(g9746)
g11249(1) = NOT(g8405)
g12036(1) = NOT(g9245)
g14110(2) = NAND(g11692, g8906)
g14741(2) = NAND(g12711, g10421)
g12879(1) = NOT(g10381)
g14892(2) = NAND(g12700, g12515)
g12878(1) = NOT(g10386)
g12337(2) = NOT(g9340)
I14650(1) = NOT(g9340)
g12886(1) = NOT(g10393)
g14758(2) = NAND(g7704, g12405)
g14226(1) = NOT(g11618)
g14683(2) = NAND(g12553, g12443)
g13889(2) = NAND(g11566, g11435)
g10572(1) = NOT(g10233)
g11534(2) = NAND(g7121, g8958)
g12972(2) = NAND(g7209, g10578)
g10877(1) = NOT(I14079)
I14705(1) = NOT(g7717)
g11404(1) = NOT(g7596)
g13291(2) = NAND(g10715, g1500)
I13805(1) = NOT(g6976)
g12598(2) = NOT(g7004)
g14376(1) = NOT(g12126)
g14807(2) = NAND(g7738, g12453)
g10869(2) = AND(g7766, g5873, g5881)
g13026(1) = NOT(g11018)
g14095(1) = NOT(g11326)
g12322(1) = NOT(I15162)
g12901(1) = NOT(g10404)
g12656(2) = NOT(g7028)
g12038(1) = NOT(I14896)
g13620(1) = NOT(g10556)
g11128(1) = NOT(g7993)
g13873(2) = NAND(g11566, g11729)
g13806(1) = NOR(g11245, g4076)
g11963(1) = NOT(g9153)
g13133(1) = NOT(g11330)
g12512(2) = NAND(g7766, g10312)
g10658(5) = NOT(I13979)
g13273(3) = NAND(g1459, g10699)
g14197(1) = NOT(g12160)
g10503(1) = NOT(g8879)
g14503(1) = NOT(g12256)
g12842(1) = NOT(g10355)
g11429(1) = NOT(g7616)
g12915(2) = NAND(g12806, g12632)
I14800(1) = NOT(g10107)
g11428(1) = NOT(g7615)
g12893(1) = NOT(g10391)
g14069(2) = NAND(g11653, g8864)
g13315(3) = NAND(g1459, g10715)
g12865(1) = NOT(g10372)
g13504(1) = NOT(g11303)
I14346(1) = NOT(g10233)
g12705(2) = NOT(g7051)
g13986(2) = NAND(g10323, g11747)
g13326(2) = NOR(g10929, g10905)
g13626(1) = NOT(g11273)
g14697(2) = NAND(g12662, g12824)
g12218(1) = NOT(I15073)
g12837(1) = NOT(g10354)
g13995(1) = NOT(g11261)
g10597(1) = NOT(g10233)
g11512(1) = NOT(g7634)
g13464(4) = NAND(g10831, g4793, g4776)
I15831(1) = NOT(g10416)
I15316(1) = NOT(g10087)
g14950(2) = NAND(g7812, g12632)
g12075(1) = NOT(I14935)
g11498(10) = NOT(I14475)
g14231(1) = NOT(g12246)
g14855(2) = NAND(g12700, g12824)
g12037(1) = NOT(I14893)
g14996(2) = NAND(g12662, g10312)
g13846(3) = NAND(g1116, g10649)
g12367(1) = NOT(I15205)
g13736(1) = NOT(g11313)
g13951(2) = NAND(g10295, g11729)
g12836(1) = NOT(g10351)
I15295(1) = NOT(g8515)
g11234(1) = NOT(g8355)
g13132(1) = NOT(g10632)
g12941(2) = NAND(g7167, g10537)
g13869(1) = NOT(g10831)
g14431(1) = NOT(g12208)
g11868(1) = NOT(g9185)
g12864(1) = NOT(g10373)
g13868(1) = NOT(g11493)
g12749(2) = NOT(g7074)
g14804(2) = NAND(g12651, g12798)
g11709(4) = NOT(I14584)
I14006(1) = NOT(g9104)
g11471(1) = NOT(g7626)
g12012(1) = NOT(g9213)
g12900(1) = NOT(g10406)
g13000(2) = NAND(g7228, g10598)
I16010(1) = NOT(g11148)
g10487(1) = NOT(g10233)
g10502(1) = NOT(g8876)
I14690(1) = NOT(g9340)
g12874(1) = NOT(g10383)
g12009(2) = NOT(I14862)
g13948(2) = NAND(g11610, g8864)
g12892(1) = NOT(g10398)
g13915(2) = NAND(g11566, g11473)
g11425(1) = NOT(g7640)
g10815(1) = NOT(g9917)
g12914(1) = NOT(g12235)
g12907(1) = NOT(g10415)
g14956(2) = NAND(g12604, g10281)
g12074(1) = NOT(I14932)
g13983(2) = NAND(g11658, g8906)
g14959(2) = NAND(g12695, g12798)
g12107(1) = NOT(g9687)
g13322(1) = NOT(g10918)
g11480(2) = NAND(g10323, g8906)
I14647(1) = NOT(g7717)
g12883(1) = NOT(g10390)
g7620(2) = NAND(I12097, I12098)
g14825(2) = NAND(g12806, g12680)
g11631(7) = NOT(g8595)
g10874(2) = AND(g7791, g6219, g6227)
g10531(1) = NOT(g8925)
g15036(2) = NAND(g12780, g12581)
g14133(2) = NAND(g11692, g11747)
g10685(9) = NOT(I13995)
g14186(1) = NOT(g11346)
g12906(1) = NOT(g10413)
g10417(1) = NOT(g7117)
g14732(2) = NAND(g12662, g12515)
g10762(12) = NOT(g8470)
g13976(1) = NOT(g11130)
g14015(2) = NAND(g11658, g11747)
g14659(2) = NAND(g12646, g12443)
I14663(1) = NOT(g9747)
g12921(1) = NOT(g12228)
g13255(1) = NOT(g10632)
g13679(1) = NOT(g10573)
g14055(2) = NAND(g11697, g11763)
g13188(1) = NOT(g10909)
g11686(4) = NOT(I14567)
g14154(2) = NAND(g11669, g8958)
g13385(7) = OR(g11967, g9479)
g7598(2) = NAND(I12075, I12076)
g10476(10) = AND(g7244, g7259, I13862)
g14947(2) = NAND(g12785, g10491)
I14687(1) = NOT(g7753)
g12013(1) = NOT(I14866)
g14275(1) = NOT(g12358)
g14237(1) = NOT(g11666)
g11470(1) = NOT(g7625)
g14101(2) = NAND(g11653, g11729)
g14024(2) = NAND(g7121, g11763)
g11467(1) = NOT(g7623)
g13595(1) = NOT(g10951)
g12882(1) = NOT(g10389)
g10475(1) = NOT(g8844)
g11170(2) = NOT(g8476)
I14016(1) = NOT(g9104)
g14999(2) = NAND(g12739, g12824)
I13759(1) = NOT(g6754)
g12026(1) = NOR(g9417, g9340)
g11401(1) = NOT(g7593)
g14755(2) = NAND(g12593, g12772)
g14927(2) = NAND(g12695, g10281)
I16898(1) = NOT(g10615)
I14708(1) = NOT(g9417)
g11560(1) = NOT(g7647)
g14209(1) = NOT(g11415)
g14208(1) = NOT(g11563)
g10607(1) = NOT(g10233)
g10530(1) = NOT(g8922)
g13665(1) = NOT(g11306)
g14723(2) = NAND(g7704, g12772)
g12692(2) = AND(g10323, g3522, g3530)
g13239(1) = NOT(g10632)
g13594(1) = NOT(g11012)
g11519(7) = NOT(g8481)
g13675(1) = NOT(g10556)
g10474(1) = NOT(g8841)
g13637(1) = NOT(g10556)
g14858(2) = NAND(g7766, g12515)
g10606(1) = NOT(g10233)
g13215(1) = NOT(g10909)
g13729(1) = NOT(g10951)
g13469(3) = NAND(g4983, g10862)
g13570(2) = OR(g9223, g11130)
g14192(1) = NOT(g11385)
g13432(3) = NAND(g4793, g10831)
g14968(2) = NAND(g12739, g10312)
g10553(1) = NOT(g8971)
g13217(3) = NAND(g4082, g10808)
I14668(1) = NOT(g7753)
g13664(1) = NOT(g11252)
g13597(2) = OR(g9247, g11149)
g11576(7) = NOT(g8542)
g14127(2) = NAND(g11653, g11435)
g11609(1) = NOT(g7660)
g12903(1) = NOT(g10411)
g11608(1) = NOT(g7659)
g10509(1) = NOT(g10233)
g12563(7) = NOT(g9864)
I14069(1) = NOT(g9104)
g14764(2) = NAND(g7738, g12798)
g12845(1) = NOT(g10358)
g12899(1) = NOT(g10407)
g14082(2) = NAND(g11697, g11537)
g12898(1) = NOT(g10405)
g13929(2) = NAND(g11669, g11763)
I14730(1) = NOT(g7717)
g12861(1) = NOT(g10367)
g14868(2) = NAND(g12755, g12680)
g14720(2) = NAND(g12593, g10266)
g13346(2) = NAND(g4854, g11012)
g14899(2) = NAND(g12744, g10421)
g14405(1) = NOT(g12170)
g11235(1) = NOT(I14301)
g14142(2) = NAND(g11715, g8958)
g12871(1) = NOT(g10378)
g12925(3) = OR(g8928, g10511)
g12181(1) = NOT(g9478)
g12735(2) = AND(g7121, g3873, g3881)
g12859(1) = NOT(g10366)
g12950(1) = NOT(g12708)
I14602(1) = NOT(g9340)
g14768(2) = NAND(g12662, g12571)
g12844(1) = NOT(g10360)
g11398(2) = NOT(I14409)
g11652(1) = NOT(g7674)
g13141(1) = NOT(g11374)
g12155(3) = NAND(g7753, g7717)
g14993(2) = NAND(g12695, g12453)
g14735(2) = NAND(g12739, g12571)
g14800(2) = NAND(g7704, g12443)
g12902(1) = NOT(g10409)
g15021(2) = NAND(g12711, g10341)
g11371(1) = NOT(g7565)
g12895(1) = NOT(g10403)
g14075(2) = NAND(g11658, g11527)
g10620(1) = NOT(g10233)
g14810(2) = NAND(g12700, g10312)
g14116(2) = NAND(g11697, g11584)
g11724(4) = NOT(I14593)
g11325(1) = NOT(g7543)
g12889(1) = NOT(g10396)
g12888(1) = NOT(g10395)
g14885(2) = NAND(g12651, g12505)
g14688(2) = NAND(g12604, g12453)
g14170(2) = NAND(g11715, g11537)
g11291(1) = NOT(g7526)
g14822(2) = NAND(g12755, g12632)
g13173(1) = NOT(g10632)
g12377(1) = NOR(g6856, g2748, g9708)
g10627(4) = NOT(I13968)
g12546(3) = NOT(g8740)
g13506(1) = NOT(g10808)
g12860(1) = NOT(g10368)
g15039(2) = NAND(g12755, g7142)
g12497(7) = NOT(g9780)
g14940(2) = NAND(g12744, g12581)
g10857(4) = NOT(g8712)
g14018(2) = NAND(g10323, g11483)
g14761(2) = NAND(g12651, g10281)
g11290(1) = NOT(I14326)
g13486(4) = NAND(g10862, g4983, g4966)
g10504(4) = NOT(g8763)
g11981(2) = NOT(I14823)
g14504(1) = NOT(g12361)
g12870(1) = NOT(g10374)
g12867(1) = NOT(g10375)
g12894(1) = NOT(g10401)
g13920(2) = NAND(g11621, g11483)
g14902(2) = NAND(g7791, g12581)
g10533(3) = NOT(g8795)
g13963(2) = NAND(g11715, g11584)
g13521(1) = NOT(g11357)
g12818(1) = NOT(g8792)
g14232(1) = NOT(g11083)
g11324(1) = NOT(g7542)
g13892(2) = NAND(g11653, g11473)
I14939(1) = NOT(g10216)
g13140(1) = NOT(g10632)
g12866(1) = NOT(g10369)
g14432(1) = NOT(g12311)
g14085(2) = NAND(g7121, g11584)
g14342(1) = NOT(g12163)
g13955(2) = NAND(g11621, g11527)
g12180(1) = NOT(g9477)
g13246(1) = NOT(g10939)
g10365(1) = NOT(g6867)
g11147(2) = NOT(g8417)
g12885(1) = NOT(g10382)
g11367(2) = NOT(I14381)
g15042(2) = NAND(g12806, g10491)
g13977(2) = NAND(g11610, g11729)
g12721(7) = NOT(g10061)
g13301(1) = NOT(g10862)
g13120(1) = NOT(g10632)
g11562(1) = NOT(g7648)
g12947(2) = NAND(g7184, g10561)
g12839(1) = NOT(g10350)
g12930(1) = NOT(g12347)
g14545(1) = NOT(g12768)
g15008(2) = NAND(g12780, g10341)
g12838(1) = NOT(g10353)
g14708(3) = AND(g74, g12369)
g14051(2) = NAND(g10323, g11527)
g12487(2) = NOT(g9340)
g10532(1) = NOT(g10233)
g14851(2) = NAND(g7738, g12505)
g11403(1) = NOT(g7595)
g11547(11) = NOT(I14505)
g13715(1) = NOT(g10573)
g12975(1) = NOT(g12752)
g12937(1) = NOT(g12419)
g7885(1) = NAND(I12270, I12271)
g13796(1) = NOR(g9158, g12527)
g14407(1) = NAND(g12008, g9807)
g13657(2) = OR(g7251, g10616)
g14643(1) = AND(g11998, g12023)
g13143(1) = NAND(g10695, g7661, g979, g1061)
I16111(1) = AND(g8691, g11409, g11381)
g13060(1) = AND(g8587, g11110)
g13411(1) = AND(g4955, g11834)
g14610(1) = AND(g1484, g10935)
g14867(1) = NOR(g10191, g12314)
g14165(1) = NOR(g8951, g11083)
I16695(1) = AND(g10207, g12523, g12463)
g14145(1) = NOR(g8945, g12259)
g14030(1) = OR(g11037, g11046)
g11111(2) = AND(g5297, g7004, g5283, g9780)
g14875(1) = AND(g1495, g10939)
g9972(1) = NAND(I13510, I13511)
g14218(1) = AND(g875, g10632)
g13384(1) = AND(g4944, g11804)
g14003(1) = NOR(g9003, g11083)
g13095(1) = OR(g11374, g1287)
g12982(1) = OR(g12220, g9968)
g14793(1) = NOR(g2988, g12228)
g14589(1) = AND(g10586, g10569)
g14588(1) = AND(g11957, g11974)
I16721(1) = AND(g10224, g12589, g12525)
g14506(2) = AND(g1430, g10755)
g13287(1) = AND(g1221, g11472)
g10733(2) = AND(g3639, g6905, g3625, g8542)
I16618(1) = AND(g10124, g12341, g12293)
g14874(1) = AND(g1099, g10909)
g14626(1) = NAND(g12232, g9852, g12159, g9715)
I16671(1) = AND(g10185, g12461, g12415)
g13994(1) = NOR(g4049, g11363)
I16143(1) = AND(g8751, g11491, g11445)
g14567(1) = AND(g10568, g10552)
g13038(1) = AND(g8509, g11034)
g14027(1) = NOR(g8734, g11363)
g14438(2) = AND(g1087, g10726)
g13288(1) = NAND(g10946, g1442)
g13077(1) = OR(g11330, g943)
g14566(1) = AND(g10566, g10551)
g12981(1) = OR(g12219, g9967)
g13300(1) = OR(g10656, g10676)
g11178(2) = AND(g6682, g7097, g6668, g10061)
g14585(1) = AND(g1141, g10905)
g7857(1) = NAND(I12241, I12242)
g14188(1) = NOR(g9162, g12259)
g10307(1) = NAND(I13730, I13731)
g13941(1) = OR(g11019, g11023)
g9528(1) = NAND(I13183, I13184)
g13959(1) = NOR(g3698, g11309)
g11123(2) = AND(g5644, g7028, g5630, g9864)
g13947(1) = NOR(g8948, g11083)
g13265(1) = AND(g9018, g11493)
g13296(1) = OR(g10626, g10657)
g14181(1) = NOR(g9083, g12259)
g13512(1) = NOR(g9077, g12527)
g13493(1) = AND(g9880, g11866)
g13035(1) = AND(g8497, g11033)
g14002(1) = NOR(g8681, g11083)
g13662(1) = OR(g10896, g10917)
g14093(1) = NOR(g8833, g11083)
g14637(1) = NAND(g12255, g9815)
g13523(1) = AND(g7046, g12246)
g14505(1) = NAND(g12073, g9961)
g13063(1) = AND(g8567, g10808)
g14613(1) = AND(g10602, g10585)
g14911(1) = NOR(g10213, g12364)
g13913(1) = NOR(g8859, g11083)
g13542(1) = AND(g10053, g11927)
g14675(1) = NAND(g12317, g9898)
g13436(1) = AND(g9721, g11811)
g12645(1) = NOR(g4467, g6961)
g13944(1) = NOR(g10262, g12259)
g10828(1) = AND(g6888, g7640)
g13155(1) = OR(g11496, g11546)
g9295(3) = NAND(I13066, I13067)
g13492(1) = AND(g9856, g11865)
g14028(1) = AND(g8673, g11797)
g14772(1) = NOR(g6044, g12252)
g13266(1) = NAND(g12440, g9920, g9843)
g14124(1) = NOR(g8830, g11083)
g7869(1) = NAND(I12252, I12253)
g14832(1) = AND(g1489, g10939)
g13728(1) = OR(g6804, g12527)
g13509(1) = AND(g9951, g11889)
g13508(1) = AND(g9927, g11888)
g14612(1) = AND(g11971, g11993)
g13047(1) = AND(g8534, g11042)
g14061(1) = AND(g8715, g11834)
g13762(1) = OR(g499, g12527)
g13627(1) = NAND(g11172, g8388)
g14767(1) = NOR(g10130, g12204)
g14122(1) = NOR(g8895, g12259)
g12924(1) = AND(g1570, g10980)
g13046(1) = AND(g6870, g11270)
g13540(1) = OR(g10822, g10827)
g14121(1) = NOR(g8891, g12259)
g13666(1) = NAND(g11190, g8441)
g14821(1) = NOR(g6390, g12314)
g13872(1) = NOR(g8745, g11083)
g11890(1) = AND(g7499, g9155)
g13081(1) = AND(g8626, g11122)
I16646(1) = AND(g10160, g12413, g12343)
g14036(1) = NOR(g8725, g11083)
g13821(1) = NAND(g11251, g8340)
g14190(1) = AND(g859, g10632)
g8069(1) = NAND(I12373, I12374)
g9258(1) = NAND(I13044, I13045)
g14816(1) = NOR(g10166, g12252)
g14126(1) = AND(g881, g10632)
g14644(1) = AND(g10610, g10605)
g14033(1) = NOR(g8808, g12259)
I16129(1) = AND(g8728, g11443, g11411)
g11185(3) = NOR(g8038, g8183, g6804)
g12644(1) = NAND(g10233, g4531)
g14433(1) = NAND(g12035, g9890)
g14343(1) = NAND(g11961, g9670)
g14202(1) = AND(g869, g10632)
g7897(1) = NAND(I12288, I12289)
g8010(1) = NAND(I12345, I12346)
g9975(1) = NAND(I13519, I13520)
g13248(1) = NAND(g9985, g12399, g9843)
g11166(2) = AND(g8363, g269, g8296, I14225)
g14163(1) = NOR(g8997, g12259)
g7803(1) = NAND(I12204, I12205)
g14572(1) = NAND(g12169, g9678)
g13080(1) = AND(g6923, g11357)
g13708(1) = NAND(g11200, g8507)
g9461(1) = NAND(I13140, I13141)
g13909(1) = NAND(g11396, g8847, g11674, g8803)
g13105(1) = NAND(g10671, g7675, g1322, g1404)
g14064(1) = NOR(g9214, g12259)
g10721(2) = AND(g3288, g6875, g3274, g8481)
g14687(1) = NOR(g5352, g12166)
g13940(1) = NAND(g11426, g8889, g11707, g8829)
g7879(1) = NAND(I12262, I12263)
g9750(1) = NAND(I13335, I13336)
g9912(1) = NAND(I13463, I13464)
g10041(1) = NAND(I13565, I13566)
g14180(1) = AND(g872, g10632)
g13660(1) = OR(g8183, g12527)
g13289(1) = OR(g10619, g10624)
g14378(1) = NAND(g11979, g9731)
g14791(1) = AND(g1146, g10909)
g13761(1) = OR(g490, g12527)
g14168(1) = AND(g887, g10632)
g11144(2) = AND(g239, g8136, g246, I14198)
g13867(1) = NAND(g11312, g8449)
g14333(1) = NAND(g12042, g12014, g11990, g11892)
g14278(1) = NOR(g562, g12259, g9217)
g14037(1) = NOR(g8748, g11083)
g9908(1) = NAND(I13453, I13454)
g13283(1) = NAND(g12440, g12399, g9843)
g14587(1) = AND(g10584, g10567)
g8238(1) = NAND(I12469, I12470)
g13525(1) = AND(g10019, g11911)
g14092(1) = NOR(g8774, g11083)
g13997(1) = OR(g11029, g11036)
g14091(1) = NOR(g8854, g12259)
g13919(1) = NOR(g3347, g11276)
g13383(1) = AND(g4765, g11797)
g14586(1) = AND(g11953, g11970)
g13294(1) = AND(g1564, g11513)
g13568(1) = NOR(g8046, g12527)
g14615(1) = AND(g10604, g10587)
g13989(1) = NOR(g8697, g11309)
g14000(1) = NOR(g8766, g12259)
g13093(1) = NAND(g10649, g7661, g979, g1061)
g11160(2) = AND(g6336, g7074, g6322, g10003)
g14182(1) = OR(g11741, g11721, g753)
g14177(1) = NAND(g11741, g11721, g753)
g9310(1) = NAND(I13078, I13079)
g14707(1) = NOR(g10143, g12259)
g13524(1) = AND(g9995, g11910)
g13699(1) = OR(g10921, g10947)
g8124(1) = NAND(I12402, I12403)
g9391(1) = NAND(I13110, I13111)
g14754(1) = NOR(g12821, g2988)
g14913(1) = AND(g1442, g10939)
g14614(1) = AND(g11975, g11997)
g14565(1) = AND(g11934, g11952)
g14641(1) = AND(g11994, g12020)
g13567(1) = AND(g10102, g11948)
g14546(1) = NAND(g12125, g9613)
g14537(1) = AND(g10550, g10529)
g14176(1) = NOR(g9044, g12259)
g12920(1) = AND(g1227, g10960)
g13349(1) = AND(g4933, g11780)
g13137(1) = NAND(g10699, g7675, g1322, g1404)
g13954(1) = NOR(g8663, g11276)
g13566(1) = AND(g7092, g12358)
g11139(2) = AND(g5990, g7051, g5976, g9935)
g13333(1) = AND(g4743, g11755)
g13623(1) = OR(g482, g12527)
g13946(1) = NOR(g8651, g11083)
g10756(2) = AND(g3990, g6928, g3976, g8595)
g14164(1) = NOR(g9000, g12259)
g14094(1) = NOR(g8770, g11083)
g12910(1) = NAND(g11002, g10601)
g14596(1) = NAND(g12196, g9775, g12124, g9663)
g13345(1) = AND(g4754, g11773)
g11025(1) = OR(g2980, g7831)
g14178(1) = NOR(g8899, g11083)
g13048(1) = AND(g8558, g11043)
g9830(1) = NAND(I13402, I13403)
g13850(1) = NAND(g11279, g8396)
g13124(1) = NAND(g10666, g7661, g979, g1061)
g14062(1) = OR(g11047, g11116)
g13507(1) = AND(g7023, g12198)
g8737(3) = NAND(I12729, I12730)
g14148(1) = AND(g884, g10632)
g14097(1) = AND(g878, g10632)
g13541(1) = AND(g7069, g12308)
g13473(1) = AND(g9797, g11841)
g14731(1) = NOR(g5698, g12204)
g13102(1) = NAND(g7523, g10759)
g13820(1) = OR(g11184, g9187, g12527)
g14253(1) = NOR(g10032, g12259, g9217)
g13281(1) = NAND(g10916, g1099)
g8359(2) = NAND(I12545, I12546)
g14090(1) = NOR(g8851, g12259)
g13491(1) = AND(g6999, g12160)
g13247(1) = AND(g8964, g11316)
g13324(1) = AND(g854, g11326)
g8873(3) = NAND(I12849, I12850)
g11032(1) = AND(g9354, g7717)
g14831(1) = AND(g1152, g10909)
g7823(1) = NAND(I12218, I12219)
g9825(1) = NAND(I13391, I13392)
g14001(1) = NOR(g739, g11083)
g14254(1) = NAND(g11968, g11933, g11951)
g7887(1) = NAND(I12278, I12279)
g14599(1) = NAND(g12207, g9739)
g12954(1) = OR(g12186, g9906)
g13059(1) = AND(g6900, g11303)
g13025(1) = AND(g8431, g11026)
g13006(1) = OR(g12284, g10034)
g13295(1) = OR(g10625, g10655)
g14726(1) = NOR(g10090, g12166)
g13176(1) = NAND(g10715, g7675, g1322, g1404)
g13632(1) = AND(g10232, g12228)
g14872(1) = NOR(g6736, g12364)
g14680(1) = AND(g12024, g12053)
g13973(1) = OR(g11024, g11028)
g11448(1) = NOR(g4191, g8790)
g8913(1) = NAND(I12877, I12878)
g14419(1) = NOR(g12152, g9546)
g14397(1) = NOR(g12120, g9416)
g14450(1) = NOR(g12195, g9598)
g14420(1) = NOR(g12153, g9490)
g14538(1) = NOR(g11973, g9828)
g14513(1) = NOR(g12222, g9754)
g14446(1) = NOR(g12190, g9644)
g7223(1) = NAND(I11878, I11879)
g7201(1) = NAND(I11865, I11866)
g14514(1) = NOR(g11959, g9760)
g14448(1) = NOR(g12192, g9699)
g14418(1) = NOR(g12151, g9594)
g14512(1) = NOR(g11955, g9753)
g14445(1) = NOR(g12188, g9693)
g14415(1) = NOR(g12147, g9590)
g11372(1) = OR(g490, g482, g8038)
g13091(1) = OR(g329, g319, g10796)
g14364(1) = NOR(g12083, g9415)
g14337(1) = NOR(g12049, g9284)
g14539(1) = NOR(g11977, g9833)
g14515(1) = NOR(g12225, g9761)
g14449(1) = NOR(g12194, g9653)
g14396(1) = NOR(g12119, g9489)
g14365(1) = NOR(g12084, g9339)
g13914(1) = OR(g8643, g11380)
g14416(1) = NOR(g12148, g9541)
g14394(1) = NOR(g12116, g9414)
g8871(1) = NAND(I12841, I12842)
g11771(1) = NOR(g8921, g4185)
g14393(1) = NOR(g12115, g9488)
g14362(1) = NOR(g12080, g9338)
g13938(1) = OR(g11213, g11191)
g14447(1) = NOR(g11938, g9698)
g14417(1) = NOR(g12149, g9648)
g14395(1) = NOR(g12118, g9542)
g14334(1) = NOR(g12044, g9337)
g14313(1) = NOR(g12016, g9250)
g14413(1) = NOR(g11914, g9638)
g14391(1) = NOR(g12112, g9585)
g14360(1) = NOR(g12078, g9484)
g13972(1) = OR(g11232, g11203)
g13794(1) = OR(g7396, g10684)
g14444(1) = NOR(g11936, g9692)
g14414(1) = NOR(g12145, g9639)
g14392(1) = NOR(g12114, g9537)
g14568(1) = NOR(g12000, g9915)
g14540(1) = NOR(g12287, g9834)
g14516(1) = NOR(g12227, g9704)
g14361(1) = NOR(g12079, g9413)
g14335(1) = NOR(g12045, g9283)
I14817(1) = NAND(g9962, I14816)
I14818(1) = NAND(g6513, I14816)
I14518(1) = NAND(g661, I14516)
g14367(8) = NOR(g9547, g12289)
I15299(1) = NAND(g10112, I15298)
I15300(1) = NAND(g1982, I15298)
I15089(1) = NAND(g2393, I15087)
I15088(1) = NAND(g9832, I15087)
g13795(1) = NAND(g11216, g401)
g14489(1) = NAND(g12126, g5084)
g12211(5) = NOR(g10099, g7097)
g14408(2) = NAND(g6069, g11924)
g11255(5) = NOR(g8623, g6928)
g12716(4) = NOR(g7812, g6555, g6549)
g13855(1) = NAND(g4944, g11804)
g13870(1) = NAND(g11773, g4732)
g13527(1) = NAND(g182, g168, g203, g12812)
g14317(2) = NAND(g5033, g11862)
g11207(5) = NOR(g3639, g6905)
g12059(5) = NOR(g9853, g7004)
g11590(1) = NAND(g6928, g3990, g4049)
g11626(4) = NOR(g7121, g3863, g3857)
g14713(2) = NOR(g12483, g9974)
I14398(2) = NAND(g8542, g3654)
g11194(5) = NOR(g3288, g6875)
g13937(1) = NOR(g8883, g4785, g11155)
I14734(1) = NAND(g9732, I14733)
I14735(1) = NAND(g5475, I14733)
g14379(2) = NAND(g5723, g11907)
g13854(1) = NAND(g4765, g11797)
I14481(1) = NAND(g10074, I14480)
I14482(1) = NAND(g655, I14480)
g13511(1) = NAND(g182, g174, g203, g12812)
g14642(2) = NOR(g12374, g9829)
I15287(2) = NAND(g10061, g6697)
I14206(1) = NAND(g3821, I14204)
I15307(1) = NAND(g10116, I15306)
I15241(2) = NAND(g10003, g6351)
g13495(1) = NAND(g1008, g11786, g7972)
I15341(1) = NAND(g10154, I15340)
g14248(2) = NOR(g6065, g10578)
g12067(5) = NOR(g5990, g7051)
I15335(1) = NAND(g2116, I15333)
g9966(2) = NAND(I13498, I13499)
g13667(2) = NAND(g3723, g11119)
g12101(5) = NOR(g6336, g7074)
g13739(2) = NAND(g11773, g11261)
I15263(1) = NAND(g10081, I15262)
I15264(1) = NAND(g2273, I15262)
g11225(5) = NOR(g3990, g6928)
g13501(2) = NOR(g3368, g11881)
g7133(1) = NAND(I11825, I11826)
I14992(1) = NAND(g9685, I14991)
I14993(1) = NAND(g6527, I14991)
g9904(2) = NAND(I13443, I13444)
I14229(1) = NAND(g979, I14228)
I14230(1) = NAND(g8055, I14228)
g9823(2) = NAND(I13383, I13384)
g13884(1) = NAND(g11797, g4727)
g11410(1) = NAND(g6875, g6895, g8696)
g11479(1) = NAND(g6875, g3288, g3347)
g12686(1) = NAND(g7097, g6682, g6736)
g12590(1) = NAND(g7097, g7110, g10229)
g12511(1) = NAND(g7028, g5644, g5698)
g12414(1) = NAND(g7028, g7041, g10165)
I14789(1) = NAND(g9891, I14788)
g12093(5) = NOR(g9924, g7028)
g12029(5) = NOR(g5644, g7028)
g12796(1) = NAND(g4467, g6961)
g13513(1) = NAND(g1351, g11815, g8002)
g13676(2) = NAND(g11834, g11283)
I14291(1) = NAND(g3835, I14289)
I15334(1) = NAND(g10152, I15333)
g13336(8) = NOR(g11330, g11011)
g12492(4) = NOR(g7704, g5170, g5164)
g13628(2) = NAND(g3372, g11107)
g14573(1) = NAND(g9506, g12249)
g14548(1) = NAND(g12208, g5774)
I15123(1) = NAND(g2102, I15121)
g11514(4) = NOR(g10295, g3161, g3155)
g12129(5) = NOR(g9992, g7051)
I15364(1) = NAND(g10182, I15363)
I15365(1) = NAND(g2675, I15363)
I13851(1) = NAND(g862, I13850)
g12558(4) = NOR(g7738, g5517, g5511)
I14766(1) = NAND(g5821, I14764)
I15130(1) = NAND(g2527, I15128)
I15193(2) = NAND(g9935, g6005)
I14258(1) = NAND(g8154, I14257)
I14259(1) = NAND(g3133, I14257)
g11571(4) = NOR(g10323, g3512, g3506)
g13971(1) = NOR(g8938, g4975, g11173)
g14712(2) = NOR(g12479, g9971)
g13727(1) = NAND(g174, g203, g168, g12812)
g13600(2) = NAND(g3021, g11039)
I15175(1) = NAND(g9977, I15174)
I14368(2) = NAND(g8481, g3303)
g11533(1) = NAND(g6905, g3639, g3698)
g11444(1) = NAND(g6905, g6918, g8733)
I15308(1) = NAND(g2407, I15306)
g13834(1) = NAND(g4754, g11773)
g13996(1) = NOR(g8938, g8822, g11173)
I15122(1) = NAND(g9910, I15121)
I14957(1) = NAND(g6181, I14955)
g13797(1) = NAND(g8102, g11273)
I14205(1) = NAND(g8508, I14204)
g12449(1) = NAND(g7004, g5297, g5352)
I14290(1) = NAND(g8282, I14289)
I14427(2) = NAND(g8595, g4005)
g12137(5) = NOR(g6682, g7097)
g14434(2) = NAND(g6415, g11945)
g12173(5) = NOR(g10050, g7074)
g14344(2) = NAND(g5377, g11885)
g14682(1) = NAND(g4933, g11780)
g11492(1) = NAND(g6928, g6941, g8756)
g12971(1) = NAND(g9024, g8977, g10664)
I14956(1) = NAND(g9620, I14955)
g14640(2) = NOR(g12371, g9824)
g12767(1) = NAND(g4467, g6961)
g13851(1) = NAND(g8224, g11360)
g13823(1) = NAND(g11313, g3774)
g13852(1) = NOR(g11320, g8347)
g14146(1) = NAND(g11020, g691)
g13480(2) = NOR(g3017, g11858)
g13378(8) = NOR(g11374, g11017)
g12002(5) = NOR(g5297, g7004)
g14521(1) = NAND(g12170, g5428)
I14855(1) = NAND(g5142, I14853)
g13634(2) = NAND(g11797, g11261)
g13709(2) = NAND(g11755, g11261)
I15213(1) = NAND(g10035, I15212)
I14714(1) = NAND(g5128, I14712)
g14752(2) = NOR(g12540, g10040)
I13852(1) = NAND(g7397, I13850)
g10754(1) = NAND(g7936, g7913, g8411)
g11238(5) = NOR(g8584, g6905)
g12342(1) = NAND(g7004, g7018, g10129)
I15105(2) = NAND(g9780, g5313)
I14885(1) = NAND(g5489, I14883)
I14854(1) = NAND(g9433, I14853)
g14120(1) = NAND(g11780, g4907)
I15003(1) = NAND(g9691, I15002)
g13779(2) = NAND(g11804, g11283)
g13945(1) = NAND(g691, g11740)
g14547(1) = NAND(g9439, g12201)
g13672(2) = NAND(g8933, g11261)
g14655(1) = NAND(g4743, g11755)
g11217(5) = NOR(g8531, g6875)
g12609(4) = NOR(g7766, g5863, g5857)
g13911(1) = NAND(g11834, g4917)
g13886(1) = NAND(g11804, g4922)
I15147(2) = NAND(g9864, g5659)
I15004(1) = NAND(g1700, I15002)
I15176(1) = NAND(g2661, I15174)
g14520(1) = NAND(g9369, g12163)
I14187(1) = NAND(g3470, I14185)
g14089(1) = NAND(g11755, g4717)
g14679(2) = NOR(g12437, g9911)
I14884(1) = NAND(g9500, I14883)
g13742(2) = NAND(g11780, g11283)
I14765(1) = NAND(g9808, I14764)
I14186(1) = NAND(g8442, I14185)
g14228(2) = NOR(g5719, g10561)
g14212(2) = NOR(g5373, g10537)
g14611(2) = NOR(g12333, g9749)
g13939(1) = NOR(g4899, g8822, g11173)
I15129(1) = NAND(g9914, I15128)
I14351(1) = NAND(g8890, I14350)
I14352(1) = NAND(g8848, I14350)
I14510(1) = NAND(g8721, I14508)
g12577(1) = NAND(g7051, g5990, g6044)
g12462(1) = NAND(g7051, g7064, g10190)
I15080(1) = NAND(g1968, I15078)
g14194(2) = NOR(g5029, g10515)
g12667(4) = NOR(g7791, g6209, g6203)
I15342(1) = NAND(g2541, I15340)
g12491(1) = NAND(g7285, g4462, g6961)
g12819(1) = NAND(g9848, g6961)
I14517(1) = NAND(g10147, I14516)
g12524(1) = NAND(g7074, g7087, g10212)
g13764(1) = NAND(g11252, g3072)
I15043(1) = NAND(g1834, I15041)
g13712(2) = NAND(g8984, g11283)
g14279(10) = NAND(g12111, g9246)
g10775(1) = NAND(g7960, g7943, g8470)
I14790(1) = NAND(g6167, I14788)
g14601(1) = NAND(g12318, g6466)
I15079(1) = NAND(g9827, I15078)
g14638(1) = NAND(g9626, g12361)
g13518(2) = NOR(g3719, g11903)
I14509(1) = NAND(g370, I14508)
I15042(1) = NAND(g9752, I15041)
I15255(1) = NAND(g1848, I15253)
I14248(1) = NAND(g1322, I14247)
I14249(1) = NAND(g8091, I14247)
g13871(1) = NAND(g4955, g11834)
g13908(1) = NOR(g4709, g8796, g11155)
g13822(1) = NAND(g8160, g11306)
g14600(1) = NAND(g9564, g12311)
I14170(1) = NAND(g8389, I14169)
I14171(1) = NAND(g3119, I14169)
I15053(1) = NAND(g2259, I15051)
I15254(1) = NAND(g10078, I15253)
g13910(1) = NOR(g4899, g4975, g11173)
g14272(2) = NOR(g6411, g10598)
I14713(1) = NAND(g9671, I14712)
I15052(1) = NAND(g9759, I15051)
I14925(1) = NAND(g5835, I14923)
g13798(1) = NAND(g11280, g3423)
g14574(1) = NAND(g12256, g6120)
I14610(1) = NAND(g8993, I14609)
I14611(1) = NAND(g8678, I14609)
I15214(1) = NAND(g1714, I15212)
g12628(1) = NAND(g7074, g6336, g6390)
I14276(1) = NAND(g8218, I14275)
I14277(1) = NAND(g3484, I14275)
g13883(1) = NOR(g4709, g4785, g11155)
g10737(1) = NAND(g6961, g9848)
I14924(1) = NAND(g9558, I14923)
g14678(2) = NOR(g12432, g9907)
g13970(1) = NOR(g8883, g8796, g11155)
g13831(1) = NOR(g11245, g7666)
g10336(1) = NAND(I13750, I13751)
g12123(1) = NOR(g6856, g2748)
g14792(1) = NOR(g10653, g10623, g10618, g10611)
g14751(1) = NOR(g10622, g10617, g10609, g10603)
g10384(1) = NOT(I13802)
g16066(2) = NOR(g10929, g13307)
g17467(1) = NOT(g14339)
g17494(1) = NOT(g14339)
I16688(1) = NOT(g10981)
I16471(1) = NOT(g12367)
g11931(1) = NOT(I14749)
g13943(1) = NOT(I16231)
g14965(2) = NAND(g12609, g12571)
g15755(1) = NOT(g13134)
g10473(1) = NOT(I13857)
g13437(20) = NOT(I15937)
g11900(2) = NOT(I14708)
g16187(2) = OR(g8822, g13486)
g17589(1) = NOT(g14981)
g17588(1) = NOT(g14782)
g17524(1) = NOT(g14933)
I15987(1) = NOT(g12381)
g14668(1) = NOT(g12450)
g11987(1) = NOT(I14833)
g17477(1) = NOT(g14848)
I15811(1) = NOT(g11128)
g11136(2) = NOT(I14192)
g14357(1) = NOT(g12181)
g14309(3) = OR(g10320, g11048)
g11966(1) = NOT(I14800)
I13906(1) = NOT(g7620)
I16663(1) = NOT(g10981)
g11855(2) = NOT(I14671)
g16629(1) = NOT(g13990)
I16150(1) = NOT(g10430)
g16472(1) = NOT(g14098)
g14255(1) = NOT(g12381)
g17642(1) = NOT(g14691)
g11894(2) = NOT(I14702)
I16535(1) = NOT(g11235)
g14238(8) = NOT(g10823)
I16526(1) = NOT(g10430)
g14065(1) = NOT(g11048)
g14912(1) = NOT(I16917)
I15682(1) = NOT(g12182)
g14219(1) = NOT(g12381)
I15590(1) = NOT(g11988)
g13070(3) = NOT(g11984)
g13584(8) = NOT(g12735)
g11986(1) = NOT(I14830)
g17476(1) = NOT(g14665)
I16077(1) = NOT(g10430)
I16102(1) = NOT(g10430)
I15636(1) = NOT(g12075)
g15727(1) = OR(g13383, g13345, g13333, g11010)
g17092(1) = NOT(g14011)
g17518(1) = NOT(g14918)
g14348(8) = NOT(g10887)
g17637(1) = NOT(g12933)
g11917(2) = NOT(I14727)
g13223(15) = NOT(I15800)
I16660(1) = NOT(g10981)
g11706(1) = NOT(I14579)
g16645(1) = NOT(g13756)
I15600(1) = NOT(g10430)
g16290(1) = NOT(g13260)
I15846(1) = NOT(g11183)
I16596(1) = NOT(g12640)
g13876(1) = NOT(g11432)
I16733(1) = NOT(g12026)
I16452(1) = NOT(g11182)
g15739(1) = NOT(g13284)
g15562(1) = NOT(g14943)
g17415(1) = NOT(g14797)
I15550(1) = NOT(g10430)
I16502(1) = NOT(g10430)
I15932(1) = NOT(g12381)
g14630(1) = NOT(g12402)
g17576(1) = NOT(g14953)
g17585(1) = NOT(g14974)
I15773(1) = NOT(g10430)
I15942(1) = NOT(g12381)
g14166(1) = NOT(g11048)
I16468(1) = NOT(g12760)
g17609(1) = NOT(g14817)
I16613(1) = NOT(g10430)
g14978(2) = NAND(g12716, g10491)
I15667(1) = NOT(g12143)
g15628(2) = NOR(g11907, g14228)
I16479(1) = NOT(g10430)
I15843(1) = NOT(g11181)
g16658(1) = NOT(g14157)
g13278(1) = NOT(g10738)
I16486(1) = NOT(g11204)
g14262(8) = NOT(g10838)
g17213(2) = NOR(g11107, g13501)
g16430(1) = OR(g182, g13657)
g16197(1) = NOT(g13861)
g13975(1) = NOT(g11048)
g16527(1) = NOT(g14048)
I16676(1) = NOT(g10588)
I15921(1) = NOT(g12381)
g10348(1) = NOT(I13762)
g15027(2) = NAND(g12667, g10341)
g11875(2) = NOT(I14687)
I15556(1) = NOT(g11928)
I17416(1) = NOT(g13806)
g12108(1) = NOT(I14964)
g17414(1) = NOT(g14627)
g14119(1) = OR(g10776, g8703)
g15995(4) = AND(g13314, g1157, g10666)
I16117(1) = NOT(g10430)
g17584(1) = NOT(g14773)
g17759(1) = NOT(g14864)
g16526(1) = NOT(g13898)
g17758(1) = NOT(g14861)
g13334(1) = NOT(g11048)
I15587(1) = NOT(g11985)
g17652(1) = NOT(g15033)
g16689(1) = NOT(g13923)
g16280(1) = NOT(g13330)
g14045(2) = NAND(g11571, g11747)
I16579(1) = NOT(g10981)
g14184(1) = NOT(g12381)
g13117(1) = NOT(g10981)
g14297(8) = NOT(g10869)
I15569(1) = NOT(g11965)
g13494(1) = NOT(g11912)
I15814(1) = NOT(g11129)
g16090(2) = NOR(g10961, g13315)
g12183(1) = NOT(I15033)
g14639(1) = NOT(I16747)
g11772(1) = NOT(I14623)
g16511(1) = NOT(g14130)
I16057(1) = NOT(g10430)
I15929(1) = NOT(g10430)
I15981(1) = NOT(g11290)
g11872(2) = NOT(I14684)
g14072(2) = NAND(g11571, g11483)
g11852(2) = NOT(I14668)
g16261(2) = OR(g7898, g13469)
g15030(2) = NAND(g12716, g12680)
g16773(1) = NOT(g14021)
g13526(1) = OR(g209, g10685, g301)
g11720(1) = NOT(I14589)
g16655(1) = NOT(g14151)
g11237(1) = NOT(I14305)
g17473(1) = NOT(g14841)
g14321(8) = NOT(g10874)
g14584(1) = NOT(g11048)
g14744(1) = NOT(g12578)
g15655(1) = NOT(g13202)
I15727(1) = NOT(g10981)
I16555(1) = NOT(g10430)
g13222(1) = NOT(g10590)
g14562(1) = NOT(g12036)
I16492(1) = NOT(g12430)
I15821(1) = NOT(g11143)
g14833(4) = NOT(g11405)
I16593(1) = NOT(g10498)
g11790(2) = NOT(I14630)
g17648(1) = NOT(g15024)
I15834(1) = NOT(g11164)
g16740(1) = NOT(g13980)
g13555(8) = NOT(g12692)
g14038(2) = NAND(g11514, g11435)
g17718(1) = NOT(g14776)
g17521(1) = NOT(g14727)
g14136(2) = NAND(g11571, g8906)
g15479(1) = NOT(g14895)
I15593(1) = NOT(g11989)
g13530(8) = NOT(g12641)
g11829(2) = NOT(I14653)
g17573(1) = NOT(g12911)
g11920(2) = NOT(I14730)
g17389(1) = NOT(g14915)
g17612(1) = NOT(g15014)
g14066(2) = NAND(g11514, g11473)
g14541(1) = NOT(g11405)
I15918(1) = NOT(g12381)
g17777(1) = NOT(g14908)
I16512(1) = NOT(g12811)
g15740(1) = NOT(g13342)
g14113(2) = NAND(g11626, g11537)
I15474(1) = NOT(g10364)
g13474(1) = NOT(g11048)
g16814(1) = NOT(g14058)
g14173(2) = NOT(g12076)
I15869(1) = NOT(g11234)
g14936(1) = OR(g10776, g8703)
g17472(1) = NOT(g14656)
I16040(1) = NOT(g10430)
g16510(1) = NOT(g14008)
g15825(3) = NOR(g7666, g13217)
g13267(3) = NOT(I15831)
g13174(1) = NOT(g10741)
I16564(1) = NOT(g10429)
g17776(1) = NOT(g14905)
g15568(1) = NOT(g14984)
g15747(1) = NOT(g13307)
g17292(3) = AND(g1075, g13093)
g13522(1) = NOT(g10981)
g16720(1) = NOT(g14234)
g16746(1) = NOT(g14258)
I15862(1) = NOT(g11215)
g16047(4) = AND(g13322, g1500, g10699)
g16684(1) = NOT(g14223)
I15702(1) = NOT(g12217)
g14191(1) = NOT(g12381)
I15564(1) = NOT(g11949)
I13889(1) = NOT(g7598)
g16523(1) = NOT(g14041)
g13062(1) = NOT(g10981)
I15872(1) = NOT(g11236)
g15746(1) = NOT(g13121)
g14107(2) = NAND(g11571, g11527)
g17738(1) = NOT(g14813)
g17645(1) = NOT(g15018)
g13087(3) = NOT(g12012)
g17194(2) = NOR(g11039, g13480)
g14078(1) = OR(g10776, g8703)
g14032(1) = NOT(g11048)
g13574(5) = NOT(I16024)
I15878(1) = NOT(g11249)
g13051(3) = NOT(g11964)
g15005(2) = NAND(g12667, g12622)
g11820(2) = NOT(I14644)
I15906(1) = NOT(g10430)
g13412(1) = NOT(g11963)
g11737(2) = OR(g8359, g8292)
I16709(1) = NOT(g10430)
g14785(1) = NOT(g12629)
g16607(1) = NOT(g13960)
g11929(1) = NOT(I14745)
I16028(1) = NOT(g12381)
g13302(1) = NOT(g12321)
g17497(1) = NOT(g14879)
g15614(1) = NOT(g14914)
g17748(3) = NAND(g562, g14708, g12323)
g14203(1) = NOT(g12381)
I16090(1) = NOT(g10430)
I16651(1) = NOT(g10542)
g15002(2) = NAND(g12609, g10312)
I15647(1) = NOT(g12109)
g13249(1) = NOT(g10590)
I16755(1) = NOT(g12377)
g16606(1) = NOT(g14110)
I16460(1) = NOT(g10430)
g17527(1) = NOT(g14741)
I15609(1) = NOT(g12013)
I15577(1) = NOT(g10430)
g17503(1) = NOT(g14892)
g11826(2) = NOT(I14650)
g14930(2) = NAND(g12609, g12515)
g13999(1) = NOT(g11048)
g17707(1) = NOT(g14758)
g17496(1) = NOT(g14683)
g16522(1) = NOT(g13889)
g13932(1) = NOT(g11534)
g17741(1) = NOT(g12972)
I15533(1) = NOT(g11867)
I15448(1) = NOT(g10877)
g11897(2) = NOT(I14705)
g15750(1) = NOT(g13291)
g13505(1) = NOT(g10981)
g10385(1) = NOT(I13805)
g17735(1) = NOT(g14807)
g16239(2) = OR(g7892, g13432)
I15620(1) = NOT(g12038)
g14888(1) = OR(g10776, g8703)
g16509(1) = NOT(g13873)
g14700(1) = NOT(g12512)
g16311(1) = NOT(g13273)
I15623(1) = NOT(g12040)
g15011(2) = NAND(g12716, g12632)
g14160(2) = NAND(g11626, g8958)
g17721(1) = NOT(g12915)
I16163(1) = NOT(g11930)
g14714(4) = NOT(g11405)
g11793(2) = NOT(I14633)
I16120(1) = NOT(g11868)
I15765(1) = NOT(g10823)
g16583(1) = NOT(g14069)
g15756(1) = NOT(g13315)
I16538(1) = NOT(g10417)
g11317(2) = NOT(I14346)
g16743(1) = NOT(g13986)
g15731(1) = NOT(g13326)
g14150(1) = NOT(g12381)
I15626(1) = NOT(g12041)
g13323(1) = NOT(g11048)
g17502(1) = NOT(g14697)
I16498(1) = NOT(g10430)
g15017(1) = OR(g10776, g8703)
g14882(2) = NAND(g12558, g12453)
g16482(1) = NOT(g13464)
g14977(1) = OR(g10776, g8703)
g17791(1) = NOT(g14950)
g17479(1) = NOT(g14855)
g17478(1) = NOT(g14996)
g16182(1) = NOT(g13846)
g14005(2) = NAND(g11514, g11729)
g16268(3) = NOR(g7913, g13121)
I15650(1) = NOT(g12110)
I15736(1) = NOT(g12322)
I16476(1) = NOT(g10430)
g16717(1) = NOT(g13951)
g12477(1) = NOT(I15295)
g17676(1) = NOT(g12941)
g17417(1) = NOT(g14804)
g17762(1) = NOT(g13000)
g11878(2) = NOT(I14690)
g16716(1) = NOT(g13948)
g16582(1) = NOT(g13915)
g13125(3) = NOR(g7863, g10762)
g13458(1) = NOT(g11048)
g14838(2) = NAND(g12492, g12405)
g17416(1) = NOT(g14956)
g13545(5) = NOT(I16010)
g16742(1) = NOT(g13983)
g17579(1) = NOT(g14959)
g14169(1) = NOT(g12381)
I16289(1) = NOT(g12107)
g13901(1) = NOT(g11480)
g10363(1) = NOT(I13779)
I16521(1) = NOT(g10430)
g11823(2) = NOT(I14647)
g15045(2) = NAND(g12716, g7142)
g11336(7) = NOT(g7620)
g17746(1) = NOT(g14825)
I15633(1) = NOT(g12074)
g17684(1) = NOT(g15036)
g14179(1) = NOT(g11048)
g16626(1) = NOT(g14133)
I16489(1) = NOT(g12793)
g17523(1) = NOT(g14732)
I15954(1) = NOT(g12381)
I16610(1) = NOT(g10981)
g16512(1) = NOT(g14015)
g12039(1) = NOT(I14899)
g11842(2) = NOT(I14660)
g17600(1) = NOT(g14659)
I15893(1) = NOT(g10430)
I15705(1) = NOT(g12218)
g14044(1) = OR(g10776, g8703)
g11705(1) = NOT(I14576)
g11845(1) = NOT(I14663)
g13189(1) = NOT(g10762)
g16529(1) = NOT(g14055)
g16528(1) = NOT(g14154)
g15831(1) = NOT(g13385)
g11294(7) = NOT(g7598)
g13065(1) = NOT(g10476)
g15582(2) = OR(g8977, g12925)
g17530(1) = NOT(g14947)
g14845(2) = NAND(g12558, g12798)
I15617(1) = NOT(g12037)
I15915(1) = NOT(g10430)
g16602(1) = NOT(g14101)
g16774(1) = NOT(g14024)
I15782(1) = NOT(g10430)
g13037(1) = NOT(g10981)
g15669(2) = NOR(g11945, g14272)
g14921(2) = NAND(g12492, g10266)
g10727(4) = NOT(I14016)
g17606(1) = NOT(g14999)
g10347(1) = NOT(I13759)
g15591(2) = NAND(g4332, g4322, g13202)
g17390(1) = NOT(g14755)
g16027(2) = NOR(g10929, g13260)
g14063(1) = NOT(g11048)
g11744(2) = NOT(I14602)
g17522(1) = NOT(g14927)
g13305(1) = NOT(g11048)
g14873(1) = NOT(I16898)
I16135(1) = NOT(g10430)
g13036(1) = NOT(g10981)
g14291(3) = NOR(g9839, g12155)
g17673(1) = NOT(g14723)
g13485(1) = NOT(g10476)
g14034(1) = NOT(g11048)
g15574(3) = AND(g4311, g13202)
g15992(2) = NOR(g10929, g13846)
g15647(2) = NOR(g11924, g14248)
I16438(1) = NOT(g11165)
g16292(3) = NOR(g7943, g13134)
g11941(2) = NOT(I14761)
g15608(2) = NOR(g11885, g14212)
g17756(1) = NOT(g14858)
g15842(1) = NOT(g13469)
g16030(1) = NOT(g13570)
g15830(1) = NOT(g13432)
g17583(1) = NOT(g14968)
g15705(1) = NOT(g13217)
g16075(1) = NOT(g13597)
g13484(1) = NOT(g10981)
g16623(1) = NOT(g14127)
g14183(1) = NOT(g12381)
g13312(1) = NOT(g11048)
g10851(4) = NOT(I14069)
g17710(1) = NOT(g14764)
g16589(1) = NOT(g14082)
g16588(1) = NOT(g13929)
g14205(1) = NOT(g12381)
g17651(1) = NOT(g14868)
g17672(1) = NOT(g14720)
g15732(1) = OR(g13411, g13384, g13349, g11016)
g16305(1) = NOT(g13346)
g14387(3) = OR(g9086, g11048)
g17505(1) = NOT(g14899)
g14937(2) = NAND(g12667, g10421)
g16630(1) = NOT(g14142)
g13414(1) = NOT(g11048)
g17811(1) = NOT(g12925)
g13082(1) = NOT(g10981)
g13107(1) = NOT(g10476)
g17582(1) = NOT(g14768)
g14198(2) = NOT(g12180)
g10710(4) = NOT(I14006)
g14204(1) = NOT(g12155)
g17603(1) = NOT(g14993)
g14971(2) = NAND(g12667, g12581)
g17681(1) = NOT(g14735)
g18061(1) = NOT(g14800)
g14104(2) = NAND(g11514, g8864)
g17239(2) = NOR(g11119, g13518)
g17504(1) = NOT(g15021)
g13106(1) = NOT(g10981)
g13463(1) = NOT(g10476)
g16585(1) = NOT(g14075)
g14149(1) = NOT(g12381)
g17737(1) = NOT(g14810)
g16608(1) = NOT(g14116)
g12490(1) = NOT(I15316)
g15585(2) = NOR(g11862, g14194)
I15788(1) = NOT(g10430)
g17499(1) = NOT(g14885)
g17498(1) = NOT(g14688)
g16692(1) = NOT(g14170)
g17611(1) = NOT(g14822)
g13110(3) = NOR(g7841, g10741)
g17529(1) = NOT(g15039)
g17528(1) = NOT(g14940)
g16771(1) = NOT(g14018)
g17709(1) = NOT(g14761)
g16515(1) = NOT(g13486)
g14962(2) = NAND(g12558, g10281)
g16584(1) = NOT(g13920)
g17774(1) = NOT(g14902)
g16725(1) = NOT(g13963)
g16044(2) = NOR(g10961, g13861)
g16652(1) = NOT(g13892)
g14794(2) = NAND(g12492, g12772)
g14844(1) = OR(g10776, g8703)
g10499(1) = NOT(I13872)
g13061(1) = NOT(g10981)
g14889(2) = NAND(g12609, g12824)
g17144(1) = NOT(g14085)
g12077(1) = NOT(I14939)
g16605(1) = NOT(g13955)
g14139(2) = NAND(g11626, g11584)
g14876(2) = NAND(g12492, g12443)
g16072(2) = NOR(g10961, g13273)
g17687(1) = NOT(g15042)
g16473(1) = NOT(g13977)
g14079(2) = NAND(g11626, g11763)
g14924(2) = NAND(g12558, g12505)
g16173(2) = OR(g8796, g13464)
g17713(1) = NOT(g12947)
g17610(1) = NOT(g15008)
g17189(1) = NOT(g14708)
g17124(1) = NOT(g14051)
g15344(1) = NOT(g14851)
g17617(1) = AND(g7885, g13326)
g12224(1) = NAND(I15088, I15089)
g13671(1) = AND(g4498, g10532)
g16052(1) = OR(g13060, g10724)
g14988(4) = NOR(g10816, g10812, g10805)
g15106(1) = NOR(g12872, g10430)
g17418(1) = AND(g9618, g14407)
g16612(1) = AND(g5603, g14927)
g16324(1) = AND(g13657, g182)
g16534(1) = AND(g5575, g14665)
g11224(1) = NAND(I14290, I14291)
g15794(1) = AND(g3239, g14008)
g13497(1) = AND(g2724, g12155)
g17321(2) = AND(g1418, g13105)
g13032(1) = NOR(g7577, g10762)
g17401(2) = AND(g1083, g13143)
g12953(1) = AND(g411, g11048)
g17119(1) = AND(g5272, g14800)
g16766(1) = AND(g6649, g12915)
g12539(1) = NAND(I15341, I15342)
g16871(1) = AND(g6597, g14908)
g17137(1) = NAND(g13727, g13511, g13527)
g15861(1) = AND(g3957, g14170)
g15170(1) = NOR(g7118, g14279)
g17177(1) = AND(g6657, g14984)
g16591(1) = AND(g5256, g14879)
g17174(1) = NOR(g9194, g14279)
g17693(1) = AND(g1306, g13291)
g16867(1) = OR(g13493, g11045)
g15871(1) = AND(g3203, g13951)
g16800(1) = OR(g13436, g11027)
g16844(1) = AND(g7212, g13000)
g15859(1) = AND(g3610, g13923)
g13056(1) = NOR(g7400, g10741)
g15968(1) = OR(g13038, g10677)
g12851(1) = NOR(g6846, g10430)
g16699(1) = AND(g7134, g12933)
g15738(1) = AND(g1111, g13260)
g17138(1) = AND(g255, g13239)
g17682(1) = AND(g9742, g14637)
g15699(1) = AND(g1437, g13861)
g16671(1) = AND(g6275, g14817)
g16260(1) = NAND(g4888, g13910, g12088)
g13942(1) = AND(g5897, g12512)
g13156(16) = AND(g10816, g10812, g10805)
g16190(1) = AND(g14626, g11810)
g13888(1) = OR(g2941, g11691)
g14555(1) = AND(g12521, g12356, g12307, I16671)
g11962(1) = NAND(I14789, I14790)
g16211(1) = AND(g5445, g14215)
g15784(1) = AND(g3235, g13977)
g17692(1) = AND(g1124, g13307)
g13306(1) = AND(g441, g11048)
g12286(1) = NAND(I15129, I15130)
g14035(1) = AND(g699, g11048)
g12853(1) = NOR(g6848, g10430)
g16870(1) = AND(g6625, g14905)
g15700(1) = AND(g3089, g13483)
g15578(1) = NOR(g7216, g14279)
g17771(1) = AND(g13288, g13190)
g16707(1) = AND(g6641, g15033)
g16202(1) = AND(g86, g14197)
g17307(1) = AND(g9498, g14343)
g16590(1) = AND(g5236, g14683)
g16986(1) = AND(g246, g13142)
g15870(1) = AND(g3231, g13948)
g13321(1) = AND(g847, g11048)
g17574(1) = AND(g9554, g14546)
g11135(1) = NAND(I14186, I14187)
g12285(1) = NAND(I15122, I15123)
g15707(1) = AND(g4082, g13506)
g15819(1) = AND(g3251, g14101)
g15818(1) = AND(g3941, g14082)
g12100(1) = NAND(I14956, I14957)
g14608(1) = AND(g12638, g12476, g12429, I16721)
g16706(1) = AND(g6621, g14868)
g16597(1) = AND(g6263, g15021)
g15965(1) = OR(g13035, g10675)
g10472(1) = NAND(I13851, I13852)
g16885(1) = AND(g6605, g14950)
g13807(1) = AND(g4504, g10606)
g13974(1) = AND(g6243, g12578)
g12431(1) = NAND(I15254, I15255)
g16596(1) = AND(g5941, g14892)
g16243(1) = AND(g6483, g14275)
g17954(1) = NOR(g832, g14279)
g15508(1) = NOR(g10320, g14279)
g16670(1) = AND(g5953, g14999)
g16734(1) = AND(g5961, g14735)
g16930(1) = AND(g239, g13132)
g13771(1) = AND(g11441, g11355, g11302, I16111)
g16667(1) = AND(g5268, g14659)
g16965(1) = AND(g269, g13140)
g16076(1) = OR(g13081, g10736)
g15570(1) = NOR(g822, g14279)
g16619(1) = AND(g6629, g14947)
g13004(1) = NOR(g7933, g10741)
g16618(1) = AND(g6609, g15039)
g16621(1) = AND(g8278, g13821)
g17134(1) = AND(g5619, g14851)
g15839(1) = AND(g3929, g13990)
g17506(1) = AND(g9744, g14505)
g15838(1) = AND(g3602, g14133)
g12136(1) = NAND(I14992, I14993)
g11761(1) = NAND(I14610, I14611)
g15815(1) = AND(g3594, g14075)
g16531(1) = AND(g5232, g14656)
g11944(1) = NAND(I14765, I14766)
g17719(1) = AND(g9818, g14675)
g13320(1) = AND(g417, g11048)
g13094(1) = NOR(g7487, g10762)
g12028(1) = NAND(I14884, I14885)
g16639(1) = AND(g6291, g14974)
g16638(1) = AND(g6271, g14773)
g16841(1) = AND(g5913, g14858)
g11118(1) = NAND(I14170, I14171)
g13341(1) = NOR(g7863, g10762)
g15814(1) = AND(g3574, g13920)
g15807(1) = AND(g3570, g13898)
g12852(1) = NOR(g6847, g10430)
g15841(1) = AND(g4273, g13868)
g11561(1) = NAND(I14517, I14518)
g11511(1) = NAND(I14481, I14482)
g16517(1) = AND(g5248, g14797)
g14719(1) = AND(g4392, g10830)
g13564(1) = AND(g4480, g12820)
g17412(1) = NAND(g14520, g14489)
g13005(1) = NOR(g7939, g10762)
g12847(1) = NOR(g6838, g10430)
g17146(1) = AND(g5965, g14895)
g12848(1) = NOR(g6839, g10430)
g13912(1) = AND(g5551, g12450)
g16321(1) = NAND(g4955, g13996, g12088)
g16304(1) = NAND(g4765, g13970, g12054)
g16516(1) = AND(g5228, g14627)
g16422(1) = AND(g8216, g13627)
g13044(1) = NOR(g7349, g10762)
g16208(1) = AND(g3965, g14085)
g17784(1) = AND(g1152, g13215)
g16614(1) = AND(g5945, g14933)
g16970(1) = OR(g13567, g11163)
g15821(1) = AND(g3598, g14110)
g16593(1) = AND(g5599, g14885)
g13020(1) = AND(g401, g11048)
g12592(1) = NAND(I15364, I15365)
g16641(1) = AND(g6613, g14782)
g13282(1) = AND(g3546, g11480)
g12846(1) = NOR(g6837, g10430)
g16635(1) = AND(g5607, g14959)
g14511(1) = OR(g10685, g546)
g16653(1) = AND(g8343, g13850)
g15913(1) = AND(g3933, g14021)
g16474(1) = AND(g8280, g13666)
g16537(1) = AND(g5937, g14855)
g16303(1) = AND(g4527, g12921)
g13778(1) = AND(g4540, g10597)
g13998(1) = AND(g6589, g12629)
g12191(1) = NAND(I15052, I15053)
g13969(1) = OR(g11448, g8913)
g16483(1) = AND(g5224, g14915)
g16536(1) = AND(g5917, g14996)
g16702(1) = AND(g5615, g14691)
g15796(1) = AND(g3586, g14015)
g17643(1) = AND(g9681, g14599)
g15840(1) = AND(g3949, g14142)
g16673(1) = AND(g6617, g14822)
g13114(1) = NOR(g7528, g10741)
g16634(1) = AND(g5264, g14953)
g16282(1) = NAND(g4933, g13939, g12088)
g13805(1) = AND(g11489, g11394, g11356, I16129)
g16690(1) = AND(g8399, g13867)
g16592(1) = AND(g5579, g14688)
g13335(1) = NOR(g7851, g10741)
g17391(1) = AND(g9556, g14378)
g15851(1) = AND(g3953, g14157)
g15872(1) = AND(g9095, g14234)
g12144(1) = NAND(I15003, I15004)
g16507(1) = NAND(g13797, g13764)
g17500(1) = NAND(g14573, g14548)
g16731(1) = AND(g7153, g12941)
g17480(1) = AND(g9683, g14433)
g16021(1) = OR(g13047, g10706)
g16866(1) = OR(g13492, g11044)
g12336(1) = NAND(I15175, I15176)
g15912(1) = AND(g3562, g14018)
g14581(1) = AND(g12587, g12428, g12357, I16695)
g14496(1) = AND(g12411, g12244, g12197, I16618)
g17156(1) = AND(g305, g13385)
g17655(1) = AND(g7897, g13342)
g15820(1) = AND(g3578, g13955)
g12939(1) = AND(g405, g11048)
g13299(1) = AND(g437, g11048)
g16803(1) = AND(g5933, g14810)
g12066(1) = NAND(I14924, I14925)
g17469(1) = AND(g4076, g13217)
g13737(1) = AND(g4501, g10571)
g13697(1) = AND(g11166, g8608)
g17601(1) = AND(g9616, g14572)
g15881(1) = AND(g3582, g13983)
g12856(1) = NOR(g10430, g6855)
g16233(1) = AND(g6137, g14251)
g16672(1) = AND(g6295, g15008)
g16306(1) = NAND(g4944, g13971, g12088)
g13461(1) = AND(g2719, g11819)
g16513(1) = AND(g8345, g13708)
g13887(1) = AND(g5204, g12402)
g15779(1) = AND(g13909, g11214)
g13393(1) = AND(g703, g11048)
g15786(1) = AND(g13940, g11233)
g14528(1) = AND(g12459, g12306, g12245, I16646)
g17654(1) = AND(g962, g13284)
g10589(1) = OR(g7223, g7201)
g11323(1) = NAND(I14351, I14352)
g17525(1) = NAND(g14600, g14574)
g15372(1) = NOR(g817, g14279)
g17586(1) = NAND(g14638, g14601)
g14210(1) = AND(g4392, g10590)
g16896(1) = AND(g262, g13120)
g16281(1) = NAND(g4754, g13937, g12054)
g17123(1) = AND(g225, g13209)
g15803(1) = OR(g12924, g10528)
g15850(1) = AND(g3606, g14151)
g16802(1) = AND(g5567, g14807)
g16730(1) = AND(g5212, g14723)
g13656(1) = AND(g278, g11144)
g16245(1) = AND(g14278, g14708)
g14654(1) = AND(g7178, g10476)
g15594(1) = NOR(g10614, g13026, g7285)
g15793(1) = AND(g3219, g13873)
g17190(1) = NOR(g723, g14279)
g16737(1) = AND(g6645, g15042)
g14216(1) = AND(g7631, g10608)
g10543(1) = AND(g8238, g437)
g11923(1) = NAND(I14734, I14735)
g12858(1) = NOR(g10365, g10430)
g11559(1) = NAND(I14509, I14510)
g16611(1) = AND(g5583, g14727)
g13830(1) = AND(g11543, g11424, g11395, I16143)
g15856(1) = AND(g9056, g14223)
g15880(1) = AND(g3211, g13980)
g13042(1) = AND(g433, g11048)
g16199(1) = AND(g3614, g14051)
g16736(1) = AND(g6303, g15036)
g12854(1) = NOR(g6849, g10430)
g12980(1) = NOR(g7909, g10741)
g16843(1) = AND(g6251, g14864)
g17726(1) = AND(g1467, g13315)
g16764(1) = AND(g6307, g14776)
g13030(1) = AND(g429, g11048)
g16869(1) = AND(g6259, g14902)
g16586(1) = NAND(g13851, g13823)
g12855(1) = NOR(g10430, g6854)
g12482(1) = NAND(I15307, I15308)
g17153(1) = AND(g6311, g14943)
g16839(1) = OR(g13473, g11035)
g13277(1) = AND(g3195, g11432)
g14193(1) = AND(g7178, g10590)
g13853(1) = AND(g4549, g10620)
g16598(1) = AND(g6283, g14899)
g15810(1) = AND(g3937, g14055)
g16288(1) = NOR(g13794, g417)
g16532(1) = AND(g5252, g14841)
g12187(1) = NAND(I15042, I15043)
g13313(1) = AND(g475, g11048)
g15967(1) = AND(g3913, g14058)
g15754(1) = NOR(g341, g7440, g13385)
g13808(1) = AND(g4543, g10607)
g12538(1) = NAND(I15334, I15335)
g15817(1) = AND(g3921, g13929)
g14583(1) = OR(g10685, g542)
g15783(1) = AND(g3215, g14098)
g15823(1) = AND(g3945, g14116)
g11906(1) = NAND(I14713, I14714)
g16669(1) = AND(g5611, g14993)
g16842(1) = AND(g6279, g14861)
g16610(1) = AND(g5260, g14918)
g16705(1) = AND(g6299, g15024)
g12478(1) = NAND(I15299, I15300)
g17405(2) = AND(g1422, g13137)
g13031(1) = NOR(g7301, g10741)
g16258(1) = OR(g13247, g10856)
g13415(1) = AND(g837, g11048)
g16617(1) = AND(g6287, g14940)
g15678(1) = AND(g1094, g13846)
g17769(1) = AND(g1146, g13188)
g16448(1) = OR(g13287, g10934)
g13325(1) = NOR(g7841, g10741)
g16595(1) = AND(g5921, g14697)
g15875(1) = AND(g3961, g13963)
g15837(1) = AND(g3255, g14127)
g13076(1) = NOR(g7443, g10741)
g11153(1) = NAND(I14205, I14206)
g17786(1) = AND(g1489, g13216)
g12850(1) = NOR(g10430, g6845)
g16616(1) = AND(g6267, g14741)
g16704(1) = AND(g5957, g15018)
g15822(1) = AND(g3925, g13960)
g16808(1) = AND(g6653, g14825)
g16928(1) = OR(g13525, g11127)
g16642(1) = AND(g6633, g14981)
g16238(1) = NAND(g4698, g13883, g12054)
g15749(1) = AND(g1454, g13273)
g17149(1) = AND(g232, g13255)
g16927(1) = OR(g13524, g11126)
g15704(1) = AND(g3440, g13504)
g15809(1) = AND(g3917, g14154)
g11206(1) = NAND(I14276, I14277)
g15808(1) = AND(g3590, g14048)
g12849(1) = NOR(g6840, g10430)
g16519(1) = AND(g5591, g14804)
g16176(1) = AND(g14596, g11779)
g16185(1) = AND(g3263, g14011)
g17424(2) = AND(g1426, g13176)
g16518(1) = AND(g5571, g14956)
g16022(1) = OR(g13048, g10707)
g16637(1) = AND(g5949, g14968)
g15712(1) = AND(g3791, g13521)
g15914(1) = AND(g3905, g14024)
g12001(1) = NAND(I14854, I14855)
g16729(1) = AND(g5240, g14720)
g17474(1) = NAND(g14547, g14521)
g16882(1) = OR(g13508, g11114)
g13833(1) = AND(g4546, g10613)
g11980(1) = NAND(I14817, I14818)
g17198(1) = NOR(g9282, g14279)
g13221(1) = AND(g6946, g11425)
g15883(1) = AND(g9180, g14258)
g17317(2) = AND(g1079, g13124)
g16636(1) = AND(g5929, g14768)
g17057(1) = AND(g446, g13173)
g16484(1) = AND(g5244, g14755)
g11193(1) = NAND(I14258, I14259)
g16805(1) = AND(g7187, g12972)
g13377(1) = NOR(g7873, g10762)
g16674(1) = AND(g6637, g15014)
g13078(1) = NOR(g7446, g10762)
g16761(1) = AND(g7170, g12947)
g12931(1) = AND(g392, g11048)
g17753(1) = AND(g13281, g13175)
g13029(1) = AND(g8359, g11030)
g15813(1) = AND(g3247, g14069)
g15805(1) = AND(g3243, g14041)
g14681(1) = AND(g4392, g10476)
g13013(1) = NOR(g7957, g10762)
g16259(1) = NAND(g4743, g13908, g12054)
g13604(1) = AND(g4495, g10487)
g17810(1) = AND(g1495, g13246)
g13633(1) = AND(g4567, g10509)
g16883(1) = OR(g13509, g11115)
g16759(1) = AND(g5587, g14761)
g16758(1) = AND(g5220, g14758)
g13832(1) = AND(g8880, g10612)
g12979(1) = AND(g424, g11048)
g17148(1) = NOR(g827, g14279)
g15882(1) = AND(g3554, g13986)
g14261(1) = AND(g4507, g10738)
g16804(1) = AND(g5905, g14813)
g12221(1) = NAND(I15079, I15080)
g13698(1) = NOR(g528, g12527, g11185)
g16506(1) = OR(g13294, g10966)
g16959(1) = OR(g13542, g11142)
g16221(1) = AND(g5791, g14231)
g16613(1) = AND(g5925, g14732)
g15848(1) = AND(g3259, g13892)
g15804(1) = AND(g3223, g13889)
g13129(1) = NOR(g7553, g10762)
g12370(1) = NAND(I15213, I15214)
g15792(1) = OR(g12920, g10501)
g15812(1) = AND(g3227, g13915)
g13319(1) = AND(g4076, g8812, g10658, g8757)
g12436(1) = NAND(I15263, I15264)
g16535(1) = AND(g5595, g14848)
g15795(1) = AND(g3566, g14130)
g13738(1) = AND(g8880, g10572)
g16760(1) = AND(g5559, g14764)
g13290(1) = AND(g3897, g11534)
g15910(1) = OR(g13025, g10654)
g13021(1) = NOR(g7544, g10741)
g16524(1) = NAND(g13822, g13798)
g16926(1) = OR(g14061, g11804, g11780)
I18495(1) = OR(g14539, g14515, g14449)
I18543(1) = OR(g14568, g14540, g14516)
I18492(1) = OR(g14538, g14513, g14446)
I18452(1) = OR(g14514, g14448, g14418)
g16876(1) = OR(g14028, g11773, g11755)
I18449(1) = OR(g14512, g14445, g14415)
g16811(1) = OR(g8690, g13914)
I18421(1) = OR(g14447, g14417, g14395)
g14187(2) = OR(g8871, g11771)
I18385(1) = OR(g14413, g14391, g14360)
I18417(1) = OR(g14444, g14414, g14392)
g13858(2) = OR(g209, g10685)
g13700(5) = NOR(g3288, g11615)
g17595(1) = NAND(g8616, g14367)
g13119(1) = NAND(g6625, g12211, g6715, g10061)
g13100(1) = NAND(g6581, g12137, g6692, g10061)
g14490(5) = NOR(g9853, g12598)
g14306(2) = NOR(g10060, g10887)
g14830(1) = NAND(g6605, g12211, g6723, g12721)
g17312(2) = NAND(g7297, g14248)
g13968(1) = NAND(g3913, g11255, g4031, g11631)
I15242(1) = NAND(g10003, I15241)
I15243(1) = NAND(g6351, I15241)
g17284(2) = NOR(g9253, g14317)
g17217(2) = NAND(g7239, g14194)
g13772(5) = NOR(g3990, g11702)
I18529(2) = NAND(g1811, g14640)
g14854(1) = NAND(g5555, g12093, g5654, g12563)
g14425(5) = NOR(g5644, g12656)
g13067(1) = NAND(g5240, g12059, g5331, g9780)
I18633(2) = NAND(g2504, g14713)
g16319(1) = NAND(g8224, g8170, g13736)
I17404(2) = NAND(g13378, g1472)
g14399(5) = NOR(g5297, g12598)
I14400(1) = NAND(g3654, I14398)
g13866(1) = NAND(g3239, g11194, g3321, g11519)
I18536(2) = NAND(g2236, g14642)
g13131(1) = NAND(g6243, g12101, g6377, g10003)
g17287(2) = NAND(g7262, g14228)
g17493(1) = NAND(g8659, g14367)
g17492(1) = NAND(g8655, g14367)
g13066(1) = NAND(g4430, g7178, g10590)
g13824(5) = NOR(g8623, g11702)
g13539(2) = NOR(g8594, g12735)
I15194(1) = NAND(g9935, I15193)
I15195(1) = NAND(g6005, I15193)
I14399(1) = NAND(g8542, I14398)
g15715(1) = NAND(g336, g305, g13385)
g12969(1) = NAND(g4388, g7178, g10476)
g14570(1) = NAND(g3933, g11255, g4023, g8595)
g13631(2) = NOR(g8068, g10733)
g17393(2) = NOR(g9386, g14379)
I14330(2) = NAND(g225, g9966)
g14519(1) = NAND(g3889, g11225, g4000, g8595)
g14247(2) = NOR(g9934, g10869)
g14529(5) = NOR(g6336, g12749)
g16296(2) = NAND(g9360, g13501)
g11169(1) = NAND(I14229, I14230)
I15166(2) = NAND(g9904, g9823)
g13479(1) = NAND(g12686, g12639, g12590, g12526)
g13478(1) = NAND(g12511, g12460, g12414, g12344)
g13765(5) = NOR(g8531, g11615)
g13084(1) = NAND(g5587, g12093, g5677, g9864)
g14636(1) = NAND(g5595, g12029, g5677, g12563)
I17460(2) = NAND(g13378, g1300)
g14014(1) = NAND(g3199, g11217, g3298, g11519)
g14664(1) = NAND(g5220, g12059, g5339, g12497)
g12999(1) = NAND(g4392, g10476, g4401)
I17446(2) = NAND(g13336, g956)
g17399(1) = NAND(g9626, g9574, g14535)
g14674(1) = NAND(g5941, g12067, g6023, g12614)
g14946(1) = NAND(g6247, g12173, g6346, g12672)
g14271(2) = NOR(g10002, g10874)
g16278(1) = NAND(g8102, g8057, g13664)
g13603(2) = NOR(g8009, g10721)
g15721(1) = NAND(g7564, g311, g13385)
I18625(2) = NAND(g2079, g14712)
I18680(2) = NAND(g2638, g14752)
I14370(1) = NAND(g3303, I14368)
g13516(1) = NAND(g11533, g11490, g11444, g11412)
g14522(5) = NOR(g9924, g12656)
I17494(2) = NAND(g13378, g1448)
g13109(1) = NAND(g6279, g12173, g6369, g10003)
g13799(5) = NOR(g8584, g11663)
g13108(1) = NAND(g5551, g12029, g5685, g9864)
g17220(1) = NAND(g9369, g9298, g14376)
g17246(1) = NAND(g9439, g9379, g14405)
g13500(2) = NOR(g8480, g12641)
g14437(2) = NOR(g9527, g11178)
g14123(1) = NAND(g10685, g10928)
g16275(2) = NAND(g9291, g13480)
I14211(2) = NAND(g9252, g9295)
I17923(2) = NAND(g13378, g1478)
I14497(2) = NAND(g9020, g8737)
g14320(2) = NOR(g9257, g11111)
g13040(1) = NAND(g5196, g12002, g5308, g9780)
g14898(1) = NAND(g5901, g12129, g6000, g12614)
I17883(2) = NAND(g13336, g1135)
g14497(5) = NOR(g5990, g12705)
g17290(1) = NAND(g9506, g9449, g14431)
g16316(2) = NAND(g9429, g13518)
I14369(1) = NAND(g8481, I14368)
g14569(1) = NAND(g3195, g11194, g3329, g8481)
g16476(2) = NOR(g8119, g13667)
g13928(1) = NAND(g3562, g11238, g3680, g11576)
g14227(2) = NOR(g9863, g10838)
g13670(2) = NOR(g8123, g10756)
I15288(1) = NAND(g10061, I15287)
I15289(1) = NAND(g6697, I15287)
g16757(2) = NAND(g13911, g13886, g14120, g11675)
g16299(1) = NAND(g8160, g8112, g13706)
g17315(1) = NAND(g9564, g9516, g14503)
g16663(3) = NAND(g13854, g13834, g14655, g12292)
g13897(1) = NAND(g3211, g11217, g3329, g11519)
g14347(2) = NOR(g9309, g11123)
I15149(1) = NAND(g5659, I15147)
g14054(1) = NAND(g3550, g11238, g3649, g11576)
I15148(1) = NAND(g9864, I15147)
g13097(1) = NAND(g5204, g12002, g5339, g9780)
g13104(1) = NAND(g1404, g10794)
g13907(1) = NAND(g3941, g11225, g4023, g11631)
g14088(1) = NAND(g3901, g11255, g4000, g11631)
I18587(2) = NAND(g2370, g14679)
g16728(2) = NAND(g13884, g13870, g14089, g11639)
g14625(1) = NAND(g3897, g11225, g4031, g8595)
g14987(1) = NAND(g6593, g12211, g6692, g12721)
g13050(1) = NAND(g5543, g12029, g5654, g9864)
g14211(2) = NOR(g9779, g10823)
I14530(2) = NAND(g8840, g8873)
g17596(1) = NAND(g8686, g14367)
g17243(2) = NAND(g7247, g14212)
g14549(5) = NOR(g9992, g12705)
I18485(2) = NAND(g1677, g14611)
I17474(2) = NAND(g13336, g1105)
g14590(1) = NAND(g3546, g11207, g3680, g8542)
g17225(1) = NAND(g8612, g14367)
g14575(5) = NOR(g10050, g12749)
g14706(1) = NAND(g6287, g12101, g6369, g12672)
g14696(1) = NAND(g5567, g12093, g5685, g12563)
g13499(1) = NAND(g11479, g11442, g11410, g11382)
g13498(1) = NAND(g12577, g12522, g12462, g12416)
g17363(1) = NAND(g8635, g14367)
g17420(2) = NOR(g9456, g14408)
g14411(2) = NOR(g9460, g11160)
g15710(1) = NAND(g319, g13385)
g13529(1) = NAND(g11590, g11544, g11492, g11446)
g13517(2) = NOR(g8541, g12692)
g13730(5) = NOR(g3639, g11663)
I17379(2) = NAND(g13336, g1129)
g13069(1) = NAND(g5889, g12067, g6000, g9935)
g13092(1) = NAND(g1061, g10761)
I15106(1) = NAND(g9780, I15105)
I15107(1) = NAND(g5313, I15105)
g13086(1) = NAND(g6235, g12101, g6346, g10003)
g14740(1) = NAND(g5913, g12129, g6031, g12614)
g14556(5) = NOR(g6682, g12790)
g14382(2) = NOR(g9390, g11139)
g17571(1) = NAND(g8579, g14367)
g11189(1) = NAND(I14248, I14249)
g16696(3) = NAND(g13871, g13855, g14682, g12340)
g13882(1) = NAND(g3590, g11207, g3672, g11576)
g17364(1) = NAND(g8639, g14367)
g14517(1) = NAND(g3231, g11217, g3321, g8481)
g14598(1) = NAND(g5248, g12002, g5331, g12497)
I14428(1) = NAND(g8595, I14427)
I14429(1) = NAND(g4005, I14427)
g13083(1) = NAND(g4392, g10590, g4434)
g14781(1) = NAND(g6259, g12173, g6377, g12672)
g13118(1) = NAND(g5897, g12067, g6031, g9935)
g14422(1) = NAND(g3187, g11194, g3298, g8481)
g14542(1) = NAND(g3582, g11238, g3672, g8542)
g14602(5) = NOR(g10099, g12790)
g17396(2) = NAND(g7345, g14272)
g14750(1) = NAND(g6633, g12137, g6715, g12721)
g13139(1) = NAND(g6589, g12137, g6723, g10061)
g17482(2) = NOR(g9523, g14434)
g13098(1) = NAND(g5933, g12129, g6023, g9935)
g14452(1) = NAND(g3538, g11207, g3649, g8542)
g13515(1) = NAND(g12628, g12588, g12524, g12464)
g14803(1) = NAND(g5208, g12059, g5308, g12497)
g16313(2) = NOR(g8005, g13600)
I18579(2) = NAND(g1945, g14678)
g16424(2) = NOR(g8064, g13628)
g13462(1) = NAND(g12449, g12412, g12342, g12294)
g17309(2) = NOR(g9305, g14344)
g15829(1) = NAND(g4112, g13831)
g10488(1) = NOR(g4616, g7133, g10336)
g13661(1) = NOR(g528, g11185)
g16581(1) = NOR(g13756, g8086)
g13622(1) = NOR(g278, g11166)
g12832(1) = OR(g10347, g10348)
g12833(1) = NOT(I15448)
g19408(1) = NOT(g16066)
g14454(34) = NOT(I16613)
g13543(1) = OR(g10543, g10565)
g14571(1) = NOT(I16688)
g14308(1) = NOT(I16471)
g13177(10) = NOT(I15782)
g14443(1) = NOT(I16596)
I16969(1) = NOT(g13943)
g17419(1) = NOT(g14965)
g13638(16) = NOT(I16057)
g15706(1) = AND(g13296, g13484)
g13835(10) = NOT(I16150)
I16855(1) = NOT(g10473)
g16099(1) = NOT(g13437)
g15864(2) = NAND(g14833, g12543, g12487)
g13024(1) = NOT(g11900)
g17264(3) = OR(g7118, g14309)
g20085(1) = NOT(g16187)
g20739(11) = AND(g16259, g4674)
g12301(4) = NAND(I15148, I15149)
g13250(1) = NOT(I15811)
g15844(2) = NAND(g14714, g9340, g12378)
g14424(1) = NOT(g11136)
I18063(1) = NOT(g14357)
g17616(1) = NOT(g14309)
I16590(1) = NOT(g11966)
g10544(5) = NOT(I13906)
g14544(1) = NOT(I16663)
g16162(1) = NOT(g13437)
g12983(11) = NOT(I15600)
g21250(1) = NOR(g9417, g9340, g17494)
g14383(1) = NOT(I16535)
g17733(1) = NOT(g14238)
g14358(1) = NOT(I16512)
g13605(14) = NOT(I16040)
I17744(1) = NOT(g14912)
g20751(11) = AND(g16260, g4836)
g13055(1) = NOT(I15682)
g13680(16) = NOT(I16077)
g16172(1) = NOT(g13584)
g13017(1) = NOT(I15633)
g11350(4) = NAND(I14369, I14370)
I16455(1) = NOT(g11845)
g13018(1) = NOT(I15636)
I19802(1) = NOT(g15727)
g17154(1) = NOT(g14348)
g16739(1) = NOT(g13223)
I17956(1) = NOT(g14562)
g15907(2) = NAND(g14833, g9417, g12487)
g13280(1) = NOT(I15846)
g21024(11) = AND(g16306, g4871)
g13416(14) = NOT(I15929)
g14616(8) = NOT(I16733)
g14276(1) = NOT(I16452)
g16127(1) = NOT(g13437)
g14366(1) = NOT(I16526)
I15572(1) = NOT(g10499)
g13431(1) = NOT(I15932)
g13716(10) = NOT(I16090)
g13745(10) = NOT(I16102)
g17745(1) = NOT(g14978)
g21460(1) = NOT(g15628)
g13075(1) = NOT(I15705)
g14563(1) = NOT(I16676)
I17324(1) = NOT(g14119)
g13279(1) = NOT(I15843)
I17842(1) = NOT(g13051)
g16969(1) = NOT(g14262)
g17013(1) = NOT(g14262)
g20237(1) = NOT(g17213)
g16968(1) = NOT(g14238)
g20035(1) = NOT(g16430)
g13258(1) = NOT(I15821)
g13410(1) = NOT(I15921)
g17683(1) = NOT(g15027)
g13015(1) = NOT(g11875)
g15969(8) = NOT(I17416)
g14336(1) = NOT(I16498)
g19369(1) = NOT(g15995)
g19857(2) = NAND(g13628, g16296)
g20887(11) = AND(g16282, g4864)
I16724(1) = NOT(g12108)
g13350(26) = NOT(I15906)
g12423(4) = NAND(I15242, I15243)
g12938(1) = NOT(I15556)
g16688(1) = NOT(g14045)
g19506(3) = NAND(g4087, g15825)
g17135(1) = NOT(g14297)
I17754(1) = NOT(g13494)
g14591(4) = NOT(I16709)
g19428(1) = NOT(g16090)
I18233(1) = NOT(g14639)
g13394(14) = NOT(I15915)
g13510(1) = NOT(I15981)
I18879(1) = NOT(g13267)
g20682(12) = AND(g16238, g4646)
g13014(1) = NOT(g11872)
g16721(1) = NOT(g14072)
g13007(1) = NOT(g11852)
g19533(1) = NOT(g16261)
g17507(1) = NOT(g15030)
I18148(1) = NOT(g13526)
g13041(1) = NOT(I15667)
g16180(1) = NOT(g13437)
g17789(1) = NOT(g14321)
g17121(1) = NOT(g14321)
g17268(2) = OR(g9220, g14387)
g13329(1) = NOT(I15893)
g12978(1) = NOT(I15593)
g13012(1) = NOT(I15626)
g14398(1) = NOT(I16555)
g14332(1) = NOT(I16492)
g19350(1) = AND(g15968, g13505)
g16223(1) = NOT(g13437)
g16186(1) = NOT(g13555)
I17876(1) = NOT(g13070)
g16685(1) = NOT(g14038)
g16654(1) = NOT(g14136)
g20676(2) = NAND(g14379, g17287)
g12998(1) = NOT(g11829)
g13034(1) = NOT(g11920)
g13242(3) = OR(g11336, g7601)
g12932(1) = NOT(I15550)
g16423(1) = NOT(g14066)
g13409(1) = NOT(I15918)
I16515(1) = NOT(g12477)
g16747(1) = NOT(g14113)
g13809(10) = NOT(I16135)
g16123(1) = NOT(g13530)
g13303(1) = NOT(I15869)
g14331(1) = NOT(I16489)
I17801(1) = NOT(g14936)
g16224(1) = AND(g14583, g14232)
g19364(1) = NOT(g15825)
g16579(1) = NOT(g13267)
g14330(1) = NOT(I16486)
g14315(1) = NOT(I16479)
g17147(1) = NOT(g14321)
g17754(1) = NOT(g14262)
I21162(1) = NOT(g17292)
g12946(1) = NOT(I15564)
g21163(11) = AND(g16321, g4878)
g19374(1) = NOT(g16047)
g10521(5) = NOT(I13889)
g12857(1) = NOT(I15474)
g13191(10) = NOT(I15788)
g11419(4) = NAND(I14428, I14429)
g17120(1) = NOT(g14262)
g16475(1) = NOT(g14107)
g12351(4) = NAND(I15194, I15195)
I17916(1) = NOT(g13087)
g20212(1) = NOT(g17194)
I17302(1) = NOT(g14044)
I17314(1) = NOT(g14078)
g13311(1) = NOT(I15878)
g17481(1) = NOT(g15005)
g12995(1) = NOT(g11820)
I17839(1) = NOT(g13412)
g13009(1) = NOT(I15617)
g14384(1) = NOT(I16538)
g13413(1) = NOT(g11737)
g13793(1) = NOT(I16120)
g13074(1) = NOT(I15702)
g13583(1) = NOT(I16028)
g14412(1) = NOT(I16564)
g15695(3) = NAND(g1266, g13125)
g20765(1) = NOT(g17748)
g17644(1) = NOT(g15002)
g14314(1) = NOT(I16476)
g13027(1) = NOT(I15647)
g14645(8) = NOT(I16755)
g14290(1) = NOT(I16460)
g13003(1) = NOT(I15609)
g12955(11) = NOT(I15577)
g17714(1) = NOT(g14930)
g12967(1) = NOT(g11790)
g13782(10) = NOT(I16117)
g12918(1) = NOT(I15533)
I16541(1) = NOT(g11929)
g13298(1) = NOT(I15862)
g12977(1) = NOT(I15590)
g19518(1) = NOT(g16239)
I17772(1) = NOT(g14888)
I18060(1) = NOT(g14198)
g13011(1) = NOT(I15623)
g13251(1) = NOT(I15814)
g14338(1) = NOT(I16502)
g17763(1) = NOT(g15011)
g12976(1) = NOT(I15587)
g13096(1) = NOT(I15727)
I16626(1) = NOT(g11986)
g16691(1) = NOT(g14160)
g17085(1) = NOT(g14238)
I16775(1) = NOT(g12183)
g13857(1) = NOT(I16163)
g16264(3) = NAND(g518, g9158, g13223)
g14031(1) = NOT(I16289)
g20875(11) = AND(g16281, g4681)
g16846(6) = AND(g14034, g12591, g11185)
g13144(10) = NOT(I15773)
I17834(1) = NOT(g14977)
g16769(1) = NOT(g13530)
g16768(1) = NOT(g13223)
I15494(1) = NOT(g10385)
I17873(1) = NOT(g15017)
I16160(1) = NOT(g11237)
g17815(1) = NOT(g14348)
g17677(1) = NOT(g14882)
g16651(1) = NOT(g14005)
g13271(1) = NOT(I15834)
g15962(2) = NAND(g14833, g9417, g9340)
g19407(1) = NOT(g16268)
g14307(1) = NOT(I16468)
g20734(2) = NAND(g14408, g17312)
g13101(1) = NOT(I15736)
g17772(1) = NOT(g14297)
g15811(1) = NOT(g13125)
g16310(1) = NOT(g13223)
g17638(1) = NOT(g14838)
g13010(1) = NOT(I15620)
g16958(1) = NOT(g14238)
g16096(1) = NOT(g13530)
g15877(2) = NAND(g14833, g9340, g12543)
g17014(1) = NOT(g14297)
g15853(2) = NAND(g14714, g9417, g12337)
g14363(1) = NOT(I16521)
g17720(1) = NOT(g15045)
I17733(1) = NOT(g14844)
g13023(1) = NOT(g11897)
I16544(1) = NOT(g11931)
g14423(1) = NOT(I16579)
I16679(1) = NOT(g12039)
g14543(1) = NOT(I16660)
g13016(1) = NOT(g11878)
g21277(1) = NOR(g9417, g9340, g17467)
I16629(1) = NOT(g11987)
g13460(1) = NOT(I15942)
g14442(1) = NOT(I16593)
g21306(1) = NOT(g15582)
g17122(1) = NOT(g14348)
g17641(1) = NOT(g14845)
g13138(1) = NOT(I15765)
g17136(1) = NOT(g14348)
g16171(1) = NOT(g13530)
I19762(1) = NOT(g15732)
g21556(1) = NOT(g15669)
g17575(1) = NOT(g14921)
g19614(2) = NAND(g1542, g16047)
g13477(1) = NOT(I15954)
g19071(2) = NOT(g15591)
g16159(1) = NOT(g13584)
g13022(1) = NOT(g11894)
g16158(1) = NOT(g13555)
g19355(1) = NOT(g16027)
g18088(2) = NOT(g13267)
g16680(1) = NOT(g13223)
g12940(1) = NOT(g11744)
g20871(2) = NAND(g14434, g17396)
g16966(1) = NOT(g14291)
g13064(1) = NOT(g11705)
g14453(1) = NOT(I16610)
g16289(1) = NOT(g13223)
g13008(1) = NOT(g11855)
g15867(2) = NAND(g14714, g9417, g9340)
g20645(2) = NAND(g14344, g17243)
g19146(1) = NOT(g15574)
g19738(1) = NOT(g15992)
g21510(1) = NOT(g15647)
g12951(1) = NOT(I15569)
g18935(2) = AND(g4322, g15574)
g19427(1) = NOT(g16292)
g16195(1) = NOT(g13437)
g13211(3) = OR(g11294, g7567)
g21430(1) = NOT(g15608)
g16124(1) = NOT(g13555)
g13304(1) = NOT(I15872)
I18370(1) = NOT(g14873)
g13028(1) = NOT(I15650)
g14536(1) = NOT(I16651)
g14252(1) = NOT(I16438)
I17989(1) = NOT(g14173)
g16853(1) = NOT(g13584)
g19597(2) = NAND(g1199, g15995)
g16809(1) = NOT(g14387)
g17717(1) = NOT(g14937)
g12997(1) = NOT(g11826)
g16712(1) = NOT(g13223)
g21012(11) = AND(g16304, g4688)
g19795(2) = NAND(g13600, g16275)
g12996(1) = NOT(g11823)
g17742(1) = NOT(g14971)
g12471(4) = NAND(I15288, I15289)
g16622(1) = NOT(g14104)
g17297(3) = NAND(g2729, g14291)
g20272(1) = NOT(g17239)
g13033(1) = NOT(g11917)
I18117(1) = NOT(g13302)
g15674(3) = NAND(g921, g13110)
g13514(1) = NOT(I15987)
g16200(1) = NOT(g13584)
g21413(1) = NOT(g15585)
g17056(1) = NOT(g13437)
I16698(1) = NOT(g12077)
g16214(1) = NOT(g13437)
g15799(1) = NOT(g13110)
g16646(4) = NOR(g13437, g11020, g11372)
g16235(1) = NOT(g13437)
g12968(1) = NOT(g11793)
g17087(1) = NOT(g14321)
g17602(1) = NOT(g14962)
g16206(1) = NOT(g13437)
g20619(2) = NAND(g14317, g17217)
g21389(3) = NOR(g10143, g17748, g12259)
g15833(2) = NAND(g14714, g12378, g12337)
g19751(1) = NOT(g16044)
g13045(1) = NOT(g11941)
g17599(1) = NOT(g14794)
g17086(1) = NOT(g14297)
g17680(1) = NOT(g14889)
g14753(1) = NOT(g11317)
g16812(1) = NOT(g13555)
g16514(1) = NOT(g14139)
g17308(1) = NOT(g14876)
g19362(1) = NOT(g16072)
g16724(1) = NOT(g14079)
g19875(2) = NAND(g13667, g16316)
g16325(1) = NOT(g13223)
g17392(1) = NOT(g14924)
g20070(1) = NOT(g16173)
g11389(4) = NAND(I14399, I14400)
g12239(4) = NAND(I15106, I15107)
g16633(1) = AND(g5196, g14921)
g15581(1) = NAND(g7232, g12999)
g16191(1) = AND(g5475, g14262)
I17692(1) = AND(g14988, g11450, g6756)
g17569(1) = OR(g14416, g14394, g11995, I18492)
g15903(1) = AND(g13796, g13223)
g19501(1) = OR(g16986, g14168)
g16701(1) = AND(g5547, g14845)
g16098(1) = AND(g5148, g14238)
g17488(1) = OR(g14361, g14335, g11954, I18417)
g15633(1) = AND(g3841, g13584)
g17809(1) = AND(g7873, g13125)
g15612(1) = AND(g3143, g13530)
g20131(1) = AND(g15170, g14309)
g15701(1) = AND(g3821, g13584)
g17515(3) = NOR(g13221, g10828)
g17175(1) = NOR(g1216, g13545)
g19576(1) = OR(g17138, g14202)
g15911(1) = AND(g3111, g13530)
g13019(1) = AND(g194, g11737)
g16025(1) = AND(g446, g14063)
g15785(1) = AND(g3558, g14107)
g19363(1) = OR(g17810, g14913)
g16203(1) = AND(g5821, g14297)
g15858(1) = AND(g3542, g14045)
g16226(1) = NOR(g8052, g13545)
g16427(1) = AND(g5216, g14876)
g19336(1) = OR(g17769, g14831)
g15902(1) = AND(g441, g13975)
I18620(1) = AND(g13156, g11450, g11498)
g17636(1) = AND(g10829, g13463)
g17510(1) = OR(g14393, g14362, g11972, I18449)
g15632(1) = AND(g3494, g13555)
g16287(1) = NOR(g13622, g11144)
g16024(1) = NOR(g14216, g11890)
g16520(1) = AND(g5909, g14965)
g21188(1) = AND(g7666, g15705)
g19467(1) = OR(g16896, g14097)
g16700(1) = AND(g5208, g14838)
g16126(1) = AND(g5495, g14262)
g14185(1) = AND(g8686, g11744)
g20675(1) = NAND(g14377, g17246, g9442)
g16855(1) = AND(g4392, g13107)
g15860(1) = AND(g3889, g14160)
g20733(1) = NAND(g14406, g17290, g9509)
g16801(1) = AND(g5120, g14238)
g16735(1) = AND(g6235, g15027)
I18803(1) = AND(g13156, g11450, g6756)
I18716(1) = AND(g13156, g11450, g6756)
g17625(8) = NOR(g14541, g12123)
g21285(1) = AND(g7857, g16027)
g15978(1) = AND(g246, g14032)
g15590(1) = AND(g3139, g13530)
g21011(1) = NAND(g14504, g17399, g9629)
g20187(1) = OR(g16202, g13491)
g16763(1) = AND(g6239, g14937)
I18568(1) = AND(g13156, g11450, g11498)
g14207(1) = AND(g8639, g11793)
g19874(1) = NAND(g13665, g16299, g8163)
g15876(1) = AND(g13512, g13223)
g20108(1) = AND(g15508, g11048)
I18713(1) = AND(g13156, g6767, g6756)
g14206(1) = AND(g8655, g11790)
g16237(1) = NOR(g8088, g13574)
g21333(1) = AND(g1300, g15740)
g15694(1) = AND(g457, g13437)
g17464(1) = OR(g14334, g14313, g11935, I18385)
g16884(1) = AND(g6159, g14321)
g16666(1) = AND(g5200, g14794)
I18765(1) = AND(g13156, g11450, g11498)
g14221(1) = AND(g8686, g11823)
g17770(1) = AND(g7863, g13189)
g19359(1) = OR(g17786, g14875)
g15937(1) = AND(g11950, g14387)
g16179(1) = AND(g6187, g14321)
g16178(1) = AND(g5845, g14297)
g15884(1) = AND(g3901, g14113)
g16762(1) = AND(g5901, g14930)
g15654(1) = AND(g3845, g13584)
I18762(1) = AND(g13156, g6767, g11498)
g15936(1) = AND(g475, g13999)
g19209(1) = NOR(g12971, g15614, g11320)
g16751(1) = AND(g13155, g13065)
g16807(1) = AND(g6585, g14978)
I17741(1) = AND(g14988, g11450, g11498)
g19619(1) = OR(g15712, g13080)
g17785(1) = AND(g13341, g10762)
g21332(1) = AND(g996, g15739)
g16806(1) = AND(g6247, g14971)
g21361(1) = AND(g7869, g16066)
g19903(1) = NAND(g13707, g16319, g8227)
g13252(2) = AND(g11561, g11511, g11469, g699)
g16193(1) = AND(g6533, g14348)
g16222(1) = AND(g6513, g14348)
g16703(1) = AND(g5889, g15002)
g19356(1) = OR(g17784, g14874)
g17490(1) = OR(g14364, g14337, g11958, I18421)
g15863(1) = AND(g13762, g13223)
g14220(1) = AND(g8612, g11820)
g15703(1) = AND(g452, g13437)
g17671(1) = AND(g7685, g13485)
g15935(1) = OR(g13029, g10665)
g16122(1) = AND(g9491, g14291)
g15873(1) = AND(g3550, g14072)
g15797(1) = AND(g3909, g14139)
I17606(1) = AND(g14988, g11450, g6756)
g17594(1) = OR(g14450, g14420, g12025, I18543)
g16840(1) = AND(g5467, g14262)
g19274(1) = OR(g17753, g14791)
g16192(1) = AND(g6191, g14321)
g15711(1) = AND(g460, g13437)
g15572(1) = NAND(g12969, g7219)
I18782(1) = AND(g13156, g11450, g6756)
g19344(1) = OR(g17771, g14832)
I17552(1) = AND(g13156, g11450, g11498)
g17570(1) = OR(g14419, g14397, g11999, I18495)
g15757(1) = AND(g3207, g14066)
I17542(1) = AND(g13156, g6767, g6756)
g18994(2) = OR(g16303, g13632)
g14296(1) = AND(g2638, g11897)
g15673(1) = AND(g182, g13437)
g15847(1) = AND(g3191, g14005)
g19522(1) = OR(g17057, g14180)
g16479(2) = NOR(g14719, g12490)
g17180(1) = NOR(g1559, g13574)
g16929(1) = AND(g6505, g14348)
g14257(1) = AND(g8612, g11878)
g20217(1) = OR(g16221, g13523)
g20644(1) = NAND(g14342, g17220, g9372)
g19207(1) = AND(g7803, g15992)
g14256(1) = AND(g2079, g11872)
g16204(1) = AND(g6537, g14348)
g16215(1) = NOR(g1211, g13545)
g19595(1) = OR(g17149, g14218)
g16026(1) = AND(g854, g14065)
g16212(1) = AND(g6167, g14321)
g20559(1) = AND(g336, g15831)
g21296(1) = AND(g7879, g16072)
I17575(1) = AND(g13156, g11450, g6756)
g15651(1) = AND(g429, g13414)
g15672(1) = AND(g433, g13458)
g20093(1) = AND(g15372, g14584)
I18740(1) = AND(g13156, g11450, g11498)
g20202(1) = OR(g16211, g13507)
g16765(1) = AND(g6581, g15045)
g15716(1) = AND(g468, g13437)
g19605(1) = OR(g15707, g13063)
g20870(1) = NAND(g14432, g17315, g9567)
g16128(1) = AND(g14333, g14166)
g15857(1) = AND(g3199, g14038)
g17511(1) = OR(g14396, g14365, g11976, I18452)
I18785(1) = AND(g13156, g6767, g11498)
g16810(1) = OR(g13461, g11032)
g16868(1) = AND(g5813, g14297)
g16161(1) = AND(g5841, g14297)
g15611(1) = AND(g471, g13437)
g15722(1) = AND(g464, g13437)
I17585(1) = AND(g14988, g11450, g11498)
g19856(1) = NAND(g13626, g16278, g8105)
g14222(1) = AND(g8655, g11826)
g16599(1) = AND(g6601, g15030)
g19911(1) = AND(g14707, g17748)
g16125(1) = AND(g5152, g14238)
g16023(1) = AND(g3813, g13584)
g19265(1) = NAND(g15721, g15715, g13091, g15710)
g15966(1) = AND(g3462, g13555)
g15631(1) = AND(g168, g13437)
g16668(1) = AND(g5543, g14962)
g15702(1) = NAND(g13066, g7293)
g19587(1) = OR(g15700, g13046)
g16160(1) = AND(g5499, g14262)
g21347(1) = AND(g1339, g15750)
g15679(1) = AND(g3470, g13555)
g17768(1) = AND(g13325, g10741)
I17529(1) = AND(g13156, g11450, g6756)
g19879(1) = OR(g15841, g13265)
g19488(1) = OR(g16965, g14148)
g16177(1) = AND(g5128, g14238)
g20241(1) = OR(g16233, g13541)
g15589(1) = AND(g411, g13334)
g15836(1) = AND(g3187, g14104)
g16733(1) = AND(g5893, g14889)
I18671(1) = AND(g13156, g11450, g6756)
g16485(1) = AND(g5563, g14924)
g17133(1) = AND(g10683, g13222)
g15874(1) = AND(g3893, g14079)
g15693(1) = AND(g269, g13474)
g15708(1) = NAND(g7340, g13083)
g15567(1) = AND(g392, g13312)
I18819(1) = AND(g13156, g11450, g11498)
g19557(1) = OR(g17123, g14190)
g14233(1) = AND(g8639, g11855)
g15653(1) = AND(g3119, g13530)
g16198(1) = NOR(g9247, g13574)
g15852(1) = AND(g13820, g13223)
g16184(1) = AND(g9285, g14183)
g19791(1) = AND(g14253, g17189)
g19604(1) = OR(g15704, g13059)
g16732(1) = AND(g5555, g14882)
g21302(1) = AND(g956, g15731)
g16207(1) = AND(g9839, g14204)
g15745(1) = AND(g686, g13223)
g16538(1) = AND(g6255, g15005)
g17145(1) = AND(g7469, g13249)
g17365(1) = AND(g7650, g13036)
g16183(1) = NOR(g9223, g13545)
g14316(1) = AND(g2370, g11920)
g20276(1) = OR(g16243, g13566)
g19475(1) = OR(g16930, g14126)
g19530(1) = NAND(g15829, g10841)
g17783(1) = AND(g7851, g13110)
g15849(1) = AND(g3538, g14136)
g19275(1) = AND(g7823, g16044)
g15652(1) = AND(g174, g13437)
g16227(1) = NOR(g1554, g13574)
g16163(1) = AND(g14254, g14179)
g15613(1) = AND(g3490, g13555)
g21378(1) = AND(g7887, g16090)
g17752(1) = AND(g7841, g13174)
g15507(1) = AND(g10970, g13305)
g16097(1) = NAND(g13319, g10998)
g21298(1) = AND(g7697, g15825)
g14295(1) = AND(g1811, g11894)
g16845(1) = AND(g6593, g15011)
g19525(1) = OR(g7696, g16811)
g17790(1) = NAND(g6311, g14575, g6322, g10003)
g15744(1) = NAND(g6641, g14602, g6719, g10061)
g15730(1) = NAND(g6609, g14556, g6711, g10061)
g19932(2) = NOR(g3376, g16296)
g15719(1) = NAND(g5256, g14490, g5335, g9780)
g20838(2) = NAND(g5041, g17284)
g13256(1) = NAND(g11846, g11294, g11812)
I18530(1) = NAND(g1811, I18529)
g17814(1) = NAND(g5579, g14522, g5673, g12563)
g17605(1) = NAND(g5559, g14425, g5630, g12563)
g13496(1) = NAND(g1351, g11336, g11815)
I18635(1) = NAND(g14713, I18633)
I17406(1) = NAND(g1472, I17404)
I18537(1) = NAND(g2236, I18536)
g15753(1) = NAND(g6239, g14529, g6351, g10003)
g20186(1) = NAND(g16926, g8177)
g20173(1) = NAND(g16696, g13972)
g16956(1) = NAND(g3925, g13824, g4019, g11631)
g13475(1) = NAND(g1008, g11294, g11786)
g13057(1) = NAND(g969, g11294)
g13459(1) = NAND(g7479, g11294, g11846)
g20011(2) = NAND(g3731, g16476)
I18634(1) = NAND(g2504, I18633)
g21124(2) = NAND(g5731, g17393)
I14332(1) = NAND(g9966, I14330)
g16625(1) = NAND(g3203, g13700, g3274, g11519)
I15168(1) = NAND(g9823, I15166)
g20717(2) = NOR(g5037, g17217)
g16741(1) = NAND(g3207, g13765, g3303, g11519)
g19981(2) = NOR(g3727, g16316)
I17462(1) = NAND(g1300, I17460)
g17755(1) = NAND(g5619, g14522, g5630, g9864)
g16875(1) = NAND(g3223, g13765, g3317, g11519)
g13079(1) = NAND(g1312, g11336)
g13476(1) = NAND(g7503, g11336, g11869)
g17744(1) = NAND(g6303, g14529, g6373, g12672)
I17447(1) = NAND(g13336, I17446)
g15735(1) = NAND(g5547, g14425, g5659, g9864)
g17846(1) = NAND(g6271, g14575, g6365, g12672)
g17686(1) = NAND(g6251, g14529, g6322, g12672)
g16854(1) = NAND(g3965, g13824, g3976, g8595)
g17514(1) = NAND(g3917, g13772, g4019, g8595)
g16694(1) = NAND(g3905, g13772, g3976, g11631)
g17788(1) = NAND(g5232, g14490, g5327, g12497)
g13130(1) = NAND(g1351, g11815, g11336)
g19611(1) = NAND(g1070, g1199, g15995)
I18627(1) = NAND(g14712, I18625)
g17773(1) = NAND(g5965, g14549, g5976, g9935)
g16815(1) = NAND(g3909, g13824, g4005, g11631)
g20979(2) = NAND(g5385, g17309)
I18681(1) = NAND(g2638, I18680)
g13264(1) = NAND(g11869, g11336, g11849)
I18626(1) = NAND(g2079, I18625)
g20995(2) = NOR(g5727, g17287)
I14331(1) = NAND(g225, I14330)
I17496(1) = NAND(g1448, I17494)
g16772(1) = NAND(g3558, g13799, g3654, g11576)
I17885(1) = NAND(g1135, I17883)
g15720(1) = NAND(g5917, g14497, g6019, g9935)
I18682(1) = NAND(g14752, I18680)
g13554(1) = NAND(g11336, g7582, g1351)
g17572(1) = NAND(g3598, g13799, g3676, g8542)
g17597(1) = NAND(g3191, g13700, g3303, g8481)
I17884(1) = NAND(g13336, I17883)
g15726(1) = NAND(g6263, g14529, g6365, g10003)
I20486(2) = NAND(g16696, g16757)
g17816(1) = NAND(g6657, g14602, g6668, g10061)
g16925(1) = NAND(g3574, g13799, g3668, g11576)
g16657(1) = NAND(g3554, g13730, g3625, g11576)
g16749(1) = NAND(g3957, g13772, g4027, g11631)
g16813(1) = NAND(g3614, g13799, g3625, g8542)
I18589(1) = NAND(g14679, I18587)
I18588(1) = NAND(g2370, I18587)
I20467(2) = NAND(g16663, g16728)
I17380(1) = NAND(g13336, I17379)
I17381(1) = NAND(g1129, I17379)
g17670(1) = NAND(g3893, g13772, g4005, g8595)
I14531(1) = NAND(g8840, I14530)
I17475(1) = NAND(g13336, I17474)
g17734(1) = NAND(g5272, g14490, g5283, g9780)
I18580(1) = NAND(g1945, I18579)
I18581(1) = NAND(g14678, I18579)
g17468(1) = NAND(g3215, g13700, g3317, g8481)
g17736(1) = NAND(g5563, g14522, g5659, g12563)
g17679(1) = NAND(g5611, g14425, g5681, g12563)
g15743(1) = NAND(g5893, g14497, g6005, g9935)
g21190(2) = NAND(g6077, g17420)
g20854(2) = NOR(g5381, g17243)
g13528(1) = NAND(g11294, g7549, g1008)
g15725(1) = NAND(g5603, g14522, g5681, g9864)
g15713(1) = NAND(g5571, g14425, g5673, g9864)
g15728(1) = NAND(g5200, g14399, g5313, g9780)
g16723(1) = NAND(g3606, g13730, g3676, g11576)
g15717(1) = NAND(g10754, g13092)
I18486(1) = NAND(g1677, I18485)
I18487(1) = NAND(g14611, I18485)
g15723(1) = NAND(g10775, g13104)
I18538(1) = NAND(g14642, I18536)
I14498(1) = NAND(g9020, I14497)
I14499(1) = NAND(g8737, I14497)
g17578(1) = NAND(g5212, g14399, g5283, g12497)
g17757(1) = NAND(g5909, g14549, g6005, g12614)
g17716(1) = NAND(g5957, g14497, g6027, g12614)
g16687(1) = NAND(g3255, g13700, g3325, g11519)
I17405(1) = NAND(g13378, I17404)
g19965(2) = NAND(g3380, g16424)
g15709(1) = NAND(g5224, g14399, g5327, g9780)
g13115(1) = NAND(g1008, g11786, g11294)
I14213(1) = NAND(g9295, I14211)
g15736(1) = NAND(g6295, g14575, g6373, g10003)
g17635(1) = NAND(g3542, g13730, g3654, g8542)
I17448(1) = NAND(g956, I17446)
g17708(1) = NAND(g5216, g14490, g5313, g12497)
g17640(1) = NAND(g5264, g14399, g5335, g12497)
I15167(1) = NAND(g9904, I15166)
g16770(1) = NAND(g3263, g13765, g3274, g8481)
g17775(1) = NAND(g6255, g14575, g6351, g12672)
I17925(1) = NAND(g1478, I17923)
g17872(1) = NAND(g6617, g14602, g6711, g12721)
g19632(1) = NAND(g1413, g1542, g16047)
I14212(1) = NAND(g9252, I14211)
I18531(1) = NAND(g14640, I18529)
I17924(1) = NAND(g13378, I17923)
g17820(1) = NAND(g5925, g14549, g6019, g12614)
I17461(1) = NAND(g13378, I17460)
g19916(2) = NAND(g3029, g16313)
g21253(2) = NAND(g6423, g17482)
g15729(1) = NAND(g5949, g14549, g6027, g9935)
I17495(1) = NAND(g13378, I17494)
g21140(2) = NOR(g6073, g17312)
I17476(1) = NAND(g1105, I17474)
g17647(1) = NAND(g5905, g14497, g5976, g12614)
g20163(1) = NAND(g16663, g13938)
g15782(1) = NAND(g6585, g14556, g6697, g10061)
g17513(1) = NAND(g3247, g13765, g3325, g8481)
g17723(1) = NAND(g6597, g14556, g6668, g12721)
g17495(1) = NAND(g3566, g13730, g3668, g8542)
g17765(1) = NAND(g6649, g14556, g6719, g12721)
g20172(1) = NAND(g16876, g8131)
g21206(2) = NOR(g6419, g17396)
I14532(1) = NAND(g8873, I14530)
g17598(1) = NAND(g3949, g13824, g4027, g8595)
g19887(2) = NOR(g3025, g16275)
g17792(1) = NAND(g6601, g14602, g6697, g12721)
g15718(1) = NOR(g13858, g11330)
g16220(1) = NOR(g13499, g4939)
g19778(1) = NOR(g16268, g1061)
g16232(1) = NOR(g13516, g4950)
g19793(1) = NOR(g16292, g1404)
g16231(1) = NOR(g13515, g4771)
g16201(1) = NOR(g13462, g4704)
g16210(1) = NOR(g13479, g4894)
g16242(1) = NOR(g13529, g4961)
g16209(1) = NOR(g13478, g4749)
g19853(1) = NOR(g15746, g1052)
g15724(1) = NOR(g13858, g11374)
g12970(1) = NOR(g10555, g10510, g10488)
g19873(1) = NOR(g15755, g1395)
g16219(1) = NOR(g13498, g4760)
g16488(1) = NOR(g13697, g13656)
g15048(1) = NOT(I16969)
g17781(1) = AND(g6772, g11592, g6789, I18785)
g17470(1) = NOT(g14454)
g16521(1) = NOT(g13543)
I18165(1) = NOT(g13177)
I18523(1) = NOT(g14443)
I18788(1) = NOT(g13138)
I18051(1) = NOT(g13680)
I18006(1) = NOT(g13638)
I20035(1) = NOT(g15706)
I17207(1) = NOT(g13835)
I18205(1) = NOT(g14563)
I17140(1) = NOT(g13835)
I18003(1) = NOT(g13638)
g20550(1) = NOT(g15864)
g15789(2) = OR(g10819, g13211)
g21393(1) = NOT(g17264)
g23393(1) = NOT(g20739)
g14669(3) = NOT(g12301)
g20269(1) = NOT(g15844)
g23630(8) = NAND(g20739, g11123)
g23067(8) = NAND(g20887, g10721)
I17154(1) = NOT(g13605)
g17466(1) = NOT(g12983)
g23112(8) = NAND(g21024, g10733)
g17657(4) = NOR(g14751, g12955)
I22725(1) = NOT(g21250)
I17114(1) = NOT(g14358)
I18320(1) = NOT(g13605)
g16540(36) = NOT(I17744)
g23425(1) = NOT(g20751)
I18034(1) = NOT(g13680)
I18408(1) = NOT(g13017)
g13877(3) = NOT(g11350)
g23733(8) = NAND(g20751, g11178)
g14277(1) = NOT(I16455)
g16640(1) = NOT(I17834)
g16676(1) = NOT(I17876)
g17700(4) = NOR(g14792, g12983)
g17766(1) = AND(g6772, g11592, g11640, I18762)
g16738(1) = NOT(I17956)
g20531(1) = NOT(g15907)
I18434(1) = NOT(g13782)
g23139(8) = NAND(g21163, g10756)
g16632(1) = NOT(g14454)
g23308(1) = NOT(g21024)
g17780(1) = AND(g6772, g11592, g11640, I18782)
g16661(1) = NOT(g14454)
I17507(1) = NOT(g13416)
I23099(1) = NOT(g20682)
g17727(4) = NOR(g12486, g12983)
g16533(1) = NOT(I17733)
I18252(1) = NOT(g13177)
I17121(1) = NOT(g14366)
g12952(1) = NOT(I15572)
I17173(1) = NOT(g13716)
I18101(1) = NOT(g13416)
I20499(1) = NOT(g16224)
I18238(1) = NOT(g13144)
I18872(1) = NOT(g13745)
g16594(1) = NOT(I17772)
I18574(1) = NOT(g13075)
g15824(1) = NOT(I17324)
g15050(1) = NOR(g12834, g13350)
g22761(1) = NOT(g21024)
I18135(1) = NOT(g13144)
I17491(1) = NOT(g13416)
g16644(1) = NOT(I17842)
I18350(1) = NOT(g13716)
I18313(1) = NOT(g13350)
I17633(1) = NOT(g13258)
g15806(1) = NOT(I17302)
g19455(2) = NAND(g15969, g10841, g7781)
I17612(1) = NOT(g13250)
g22654(3) = NOR(g7733, g19506)
I17098(1) = NOT(g14336)
I18071(1) = NOT(g13680)
g22759(1) = NOT(g19857)
g17663(4) = NOR(g10205, g12983)
g16695(1) = NOT(g14454)
I17228(1) = NOT(g13350)
g23285(1) = NOT(g20887)
g14609(1) = NOT(I16724)
I17420(1) = NOT(g13394)
I17456(1) = NOT(g13680)
I18482(1) = NOT(g13350)
g14745(3) = NOT(g12423)
I18248(1) = NOT(g12938)
I18089(1) = NOT(g13144)
g22406(1) = NOT(g19506)
I17355(1) = NOT(g14591)
g23699(8) = NAND(g21012, g11160)
I18810(1) = NOT(g13716)
g18091(1) = NOT(I18879)
g23382(1) = NOT(g20682)
I17675(1) = NOT(g13394)
I17374(1) = NOT(g13638)
I18104(1) = NOT(g13177)
I17699(1) = NOT(g13416)
g19495(2) = NAND(g15969, g10841, g7781)
I17125(1) = NOT(g13809)
g15800(2) = OR(g10821, g13242)
g14441(1) = NOT(I16590)
I17695(1) = NOT(g14330)
I17008(1) = NOT(g12857)
g16234(1) = AND(g6772, g6782, g11640, I17575)
g23666(8) = NAND(g20875, g11139)
g20192(1) = NOT(g17268)
I17661(1) = NOT(g13329)
I17615(1) = NOT(g13251)
I18310(1) = NOT(g12978)
g17690(1) = AND(g11547, g11592, g11640, I18671)
I18379(1) = NOT(g13012)
I17783(1) = NOT(g13304)
g16213(1) = AND(g6772, g6782, g11640, I17552)
g23909(2) = NAND(g7028, g20739)
I17181(1) = NOT(g13745)
I17671(1) = NOT(g13280)
g19063(3) = NOR(g7909, g15674)
g23949(2) = NAND(g7074, g21012)
g17491(1) = NOT(g12983)
g15816(1) = NOT(I17314)
I22024(1) = NOT(g19350)
g16580(1) = NOT(I17754)
g22845(1) = NOT(g20682)
g17794(14) = NOT(g13350)
g14676(1) = NOT(I16775)
g17694(4) = NOR(g12435, g12955)
I18323(1) = NOT(g13680)
g22718(1) = NOT(g20887)
I17094(1) = NOT(g14331)
I17658(1) = NOT(g13394)
g23400(1) = NOT(g20676)
g17653(1) = AND(g11547, g11592, g6789, I18620)
I18259(1) = NOT(g12946)
g15580(1) = NOT(g13242)
I18852(1) = NOT(g13716)
I18120(1) = NOT(g13350)
I18301(1) = NOT(g12976)
I17763(1) = NOT(g13191)
g14359(1) = NOT(I16515)
I17425(1) = NOT(g13416)
I17118(1) = NOT(g14363)
I17111(1) = NOT(g13809)
I17590(1) = NOT(g14591)
I18031(1) = NOT(g13680)
g15079(1) = AND(g2151, g12955)
I17750(1) = NOT(g14383)
I17148(1) = NOT(g14442)
g23082(1) = NOT(g21024)
I18526(1) = NOT(g13055)
I18868(1) = NOT(g14315)
g22858(1) = NOT(g20751)
g16615(1) = NOT(I17801)
g22844(1) = NOT(g21163)
I18832(1) = NOT(g13782)
g23972(2) = NAND(g7097, g20751)
g23286(2) = NAND(g6875, g20887)
I17159(1) = NOT(g13350)
I18151(1) = NOT(g13144)
g23626(2) = NOR(g17309, g20854)
g15084(1) = AND(g2710, g12983)
g17058(1) = NOT(I18148)
g17301(1) = NOT(g14454)
g13933(3) = NOT(g11419)
g23605(1) = NOT(g20739)
g16727(1) = NOT(g14454)
g14701(3) = NOT(g12351)
I18078(1) = NOT(g13350)
g20375(3) = AND(g671, g16846)
g17747(1) = AND(g6772, g11592, g11640, I18740)
g13856(1) = NOT(I16160)
I18364(1) = NOT(g13009)
g17366(1) = NOT(g14454)
I17780(1) = NOT(g13303)
I18125(1) = NOT(g13191)
g15122(1) = NOR(g6959, g13605)
g23590(8) = NAND(g20682, g11111)
g16873(1) = NOT(I18063)
g17817(1) = AND(g11547, g6782, g11640, I18819)
I17131(1) = NOT(g14384)
g14510(1) = NOT(I16629)
g16726(1) = NOT(g14454)
I18224(1) = NOT(g13793)
I18571(1) = NOT(g13074)
g16320(1) = NOT(g14454)
g16530(1) = NOT(g14454)
g20000(3) = NOR(g13661, g16264)
g23108(2) = NOR(g16424, g19932)
I17143(1) = NOT(g14412)
g19513(2) = NAND(g15969, g10841, g10922)
I18842(1) = NOT(g13809)
g19524(1) = NOT(g15695)
g15078(1) = AND(g10361, g12955)
g16283(1) = AND(g11547, g11592, g6789, I17606)
I18280(1) = NOT(g12951)
g23563(1) = NOT(g20682)
I18865(1) = NOT(g14314)
g22870(1) = NOT(g20887)
g19546(2) = NAND(g15969, g10841, g10884)
g17197(1) = NOT(I18233)
g17411(1) = NOT(g14454)
I18270(1) = NOT(g13191)
g16750(1) = NOT(g14454)
g17767(1) = AND(g6772, g11592, g6789, I18765)
g19510(2) = NAND(g15969, g10841, g10899)
g20248(16) = NAND(g17056, g14146, g14123)
I18875(1) = NOT(g13782)
I18822(1) = NOT(g13745)
g15083(1) = AND(g10362, g12983)
g14385(1) = NOT(I16541)
g14564(1) = NOT(I16679)
I17747(1) = NOT(g13298)
I18469(1) = NOT(g13809)
I17639(1) = NOT(g13350)
I17704(1) = NOT(g13144)
g21451(1) = NOT(I21162)
g16872(1) = NOT(I18060)
g21062(3) = NOR(g9547, g17297)
I17128(1) = NOT(g13835)
g17157(16) = NOT(g13350)
I17442(1) = NOT(g13638)
I18285(1) = NOT(g13638)
g19140(3) = NOR(g7939, g15695)
I17136(1) = NOT(g14398)
g15060(1) = NOR(g13350, g6814)
g16767(1) = NOT(I17989)
g23978(3) = NAND(g572, g21389, g12323)
I17188(1) = NOT(g13782)
I18177(1) = NOT(g13191)
g17793(1) = AND(g6772, g11592, g6789, I18803)
I18376(1) = NOT(g14332)
I18009(1) = NOT(g13680)
g19609(1) = NOT(g16264)
I18476(1) = NOT(g14031)
g23645(1) = NOT(g20875)
g20078(1) = NOT(g16846)
I18382(1) = NOT(g13350)
I18518(1) = NOT(g13835)
I18154(1) = NOT(g13177)
g12875(2) = NOT(I15494)
g23127(1) = NOT(g21163)
g23889(1) = NOT(g20682)
I17436(1) = NOT(g13416)
g16963(1) = NOT(I18117)
I18083(1) = NOT(g13394)
g17410(1) = NOT(g12955)
g23931(1) = NOT(g20875)
g14790(1) = NOT(I16855)
I18143(1) = NOT(g13350)
I18411(1) = NOT(g13018)
g23586(2) = NOR(g17284, g20717)
g20643(1) = NOT(g15962)
I17679(1) = NOT(g13416)
I18214(1) = NOT(g12918)
I18861(1) = NOT(g14307)
I17808(1) = NOT(g13311)
I17108(1) = NOT(g13782)
g23411(1) = NOT(g20734)
I18131(1) = NOT(g13350)
g17216(1) = NOT(g14454)
I18674(1) = NOT(g13101)
g23714(1) = NOT(g20751)
g20065(1) = NOT(g16846)
g16539(1) = AND(g11547, g6782, g6789, I17741)
g23055(1) = NOT(g20887)
g17242(1) = NOT(g14454)
g20595(1) = NOT(g15877)
g20782(1) = NOT(g15853)
g23402(1) = NOT(g20875)
I17668(1) = NOT(g13279)
I18373(1) = NOT(g13011)
g17465(1) = NOT(g12955)
I17488(1) = NOT(g13394)
I17653(1) = NOT(g14276)
g14509(1) = NOT(I16626)
g17619(4) = NOR(g10179, g12955)
I18849(1) = NOT(g14290)
I18398(1) = NOT(g13745)
I18048(1) = NOT(g13638)
I18858(1) = NOT(g13835)
g16205(1) = AND(g11547, g6782, g11640, I17542)
g23341(1) = NOT(g21163)
I18829(1) = NOT(g13350)
I18221(1) = NOT(g13605)
I22769(1) = NOT(g21277)
g16708(1) = NOT(I17916)
I17249(1) = NOT(g13605)
g19483(2) = NAND(g15969, g10841, g10922)
I18344(1) = NOT(g13003)
I18341(1) = NOT(g14308)
g19061(1) = NOT(I19762)
g22492(1) = NOT(g19614)
I18028(1) = NOT(g13638)
g23063(2) = NOR(g16313, g19887)
I17650(1) = NOT(g13271)
g23932(2) = NAND(g7051, g20875)
I17723(1) = NOT(g13177)
I19917(1) = NOT(g18088)
I17104(1) = NOT(g12932)
g23423(1) = NOT(g20871)
g16631(1) = NOT(g14454)
I18262(1) = NOT(g13857)
g23908(1) = NOT(g20739)
I18307(1) = NOT(g12977)
I17636(1) = NOT(g14252)
I18839(1) = NOT(g13716)
I17198(1) = NOT(g13809)
g20328(1) = NOT(g15867)
I18446(1) = NOT(g13028)
I18443(1) = NOT(g13027)
g23391(1) = NOT(g20645)
I17976(1) = NOT(g13638)
g16643(1) = NOT(I17839)
g22311(1) = NOT(g18935)
I17101(1) = NOT(g14338)
g15571(1) = NOT(g13211)
g17724(1) = AND(g11547, g11592, g11640, I18713)
g17725(1) = AND(g11547, g11592, g6789, I18716)
g17429(1) = NOT(I18370)
g15125(1) = OR(g10363, g13605)
g14582(1) = NOT(I16698)
g16244(1) = AND(g11547, g11592, g6789, I17585)
I18855(1) = NOT(g13745)
I18367(1) = NOT(g13010)
g17613(1) = AND(g11547, g11592, g11640, I18568)
I17401(1) = NOT(g13394)
I18265(1) = NOT(g13350)
g20033(1) = NOT(g16579)
I17392(1) = NOT(g13680)
g23342(2) = NAND(g6928, g21163)
g23662(2) = NOR(g17393, g20995)
I17471(1) = NOT(g13394)
g22449(1) = NOT(g19597)
g22897(1) = NOT(g21024)
g23309(2) = NAND(g6905, g21024)
g14386(1) = NOT(I16544)
I17166(1) = NOT(g14536)
g16194(1) = AND(g11547, g6782, g11640, I17529)
g22896(1) = NOT(g21012)
g22716(1) = NOT(g19795)
g16675(1) = NOT(I17873)
g23948(1) = NOT(g21012)
I18168(1) = NOT(g13191)
g22857(1) = NOT(g20739)
g14786(3) = NOT(g12471)
I17609(1) = NOT(g13510)
g20388(1) = NOT(g17297)
I18180(1) = NOT(g13605)
g19502(1) = NOT(g15674)
g16609(1) = NOT(g14454)
g17512(1) = NOT(g12983)
g23413(1) = NOT(g21012)
g19549(2) = NAND(g15969, g10841, g10899)
g20540(1) = NOT(g16646)
g22869(1) = NOT(g20875)
g19264(1) = NOT(I19802)
g23695(2) = NOR(g17420, g21140)
g17471(1) = NOT(g14454)
g23380(1) = NOT(g20619)
g23182(1) = NOT(g21389)
g22161(3) = AND(g13202, g19071)
g20572(1) = NOT(g15833)
I17276(1) = NOT(g13605)
g22919(1) = NOT(g21163)
g20905(3) = OR(g7216, g17264)
g23890(2) = NAND(g7004, g20682)
I18479(1) = NOT(g13041)
g23971(1) = NOT(g20751)
g23135(2) = NOR(g16476, g19981)
g22842(1) = NOT(g19875)
g23681(1) = NOT(g21012)
g17489(1) = NOT(g12955)
g19589(2) = NAND(g15969, g10841, g10884)
g13902(3) = NOT(g11389)
g16486(1) = AND(g6772, g11592, g6789, I17692)
g23729(2) = NOR(g17482, g21206)
g14631(3) = NOT(g12239)
g19337(1) = OR(g17770, g17785)
g15138(1) = NOR(g13680, g6993)
g19572(1) = OR(g17133, g14193)
g22707(1) = OR(g20559, g17156)
g15069(1) = NOR(g6828, g13416)
g18655(1) = AND(g15106, g14454)
g15101(1) = NOR(g12871, g14591)
g19267(1) = OR(g17752, g17768)
g18993(1) = AND(g11224, g16172)
g15049(1) = NOR(g13350, g6799)
g20148(1) = OR(g16128, g13393)
g15074(1) = NOR(g12845, g13416)
g22680(1) = AND(g19530, g7781)
g15162(1) = NOR(g13809, g12904)
g19536(1) = AND(g518, g16768)
g19564(1) = AND(g17175, g13976)
g15063(1) = NOR(g6818, g13394)
g15144(1) = NOR(g13716, g12890)
g19062(1) = AND(g446, g16180)
g19904(1) = OR(g17636, g14654)
g17176(1) = AND(g8616, g13008)
g19756(1) = AND(g9899, g17154)
g16957(1) = AND(g13064, g10418)
g11591(1) = NAND(I14531, I14532)
g18909(1) = AND(g16226, g13570)
g19691(1) = AND(g9614, g17085)
g18974(1) = AND(g174, g16127)
g17139(1) = AND(g8635, g12967)
g18992(1) = AND(g8341, g16171)
g23392(1) = AND(g7247, g21430)
g23424(1) = AND(g7345, g21556)
g19768(1) = AND(g2803, g15833)
g15904(2) = NAND(I17380, I17381)
g15137(1) = NOR(g6992, g13680)
g15070(1) = NOR(g6829, g13416)
g15103(1) = AND(g4180, g14454)
g16119(2) = NAND(I17475, I17476)
g19717(1) = AND(g6527, g17122)
g20193(1) = AND(g15578, g17264)
g15065(1) = NOR(g13394, g12840)
g20165(1) = AND(g5156, g17733)
g16681(2) = NAND(I17884, I17885)
g15168(1) = NOR(g13835, g12909)
g17592(1) = NAND(I18530, I18531)
g23401(1) = AND(g7262, g21460)
g15089(1) = NOR(g13144, g12861)
g21276(1) = AND(g10157, g17625)
g19716(1) = AND(g12100, g17121)
g15111(1) = AND(g4281, g14454)
g19449(1) = OR(g15567, g12939)
g15052(1) = NOR(g12835, g13350)
g23900(1) = AND(g1129, g19408)
g19681(1) = AND(g5835, g17014)
g20196(1) = OR(g16207, g13497)
g15136(1) = NOR(g13680, g12885)
g15077(1) = AND(g2138, g12955)
g15145(1) = NOR(g12891, g13716)
g18982(1) = AND(g3835, g16159)
g21382(1) = AND(g10086, g17625)
g20109(1) = AND(g17954, g17616)
g17662(1) = NAND(I18634, I18635)
g20174(1) = AND(g5503, g17754)
g18949(1) = AND(g10183, g17625)
g15133(1) = NOR(g12883, g13638)
g21348(1) = AND(g10121, g17625)
g15076(1) = AND(g2130, g12955)
g16279(1) = AND(g4512, g14424)
g22760(1) = AND(g9360, g20237)
g18933(1) = AND(g16237, g13597)
g22983(1) = NOR(g979, g16268, g19853)
g20077(1) = OR(g16025, g13320)
g19461(1) = AND(g11708, g16846)
g19145(1) = AND(g8450, g16200)
g19516(1) = AND(g7824, g16097)
g19736(1) = AND(g12136, g17136)
g19393(1) = AND(g691, g16325)
g20160(1) = OR(g16163, g13415)
g15166(1) = NOR(g13835, g7096)
g19486(1) = OR(g15589, g12979)
g19555(1) = OR(g15672, g13030)
g15140(1) = NOR(g12887, g13680)
g22191(1) = AND(g8119, g19875)
g19069(1) = AND(g8397, g16186)
g17191(1) = AND(g1384, g13242)
g11545(1) = NAND(I14498, I14499)
g22534(1) = AND(g8766, g21389)
g15158(1) = NOR(g13782, g12901)
g19545(1) = AND(g3147, g16769)
g15110(1) = AND(g4245, g14454)
g15151(1) = NOR(g13745, g7027)
g17140(1) = AND(g8616, g12968)
g15161(1) = NOR(g13809, g7073)
g22871(1) = AND(g9523, g20871)
g22152(1) = OR(g21188, g17469)
g19656(1) = AND(g2807, g15844)
g23574(1) = OR(g20093, g20108)
g19680(1) = AND(g12028, g17013)
g15126(1) = NOR(g12878, g13605)
g15124(1) = OR(g13605, g4581)
g21289(1) = NAND(g14616, g17493)
g18890(1) = AND(g10158, g17625)
g15067(1) = NOR(g12842, g13394)
g15135(1) = NOR(g6990, g13638)
g16093(2) = NAND(I17461, I17462)
g15117(1) = AND(g4300, g14454)
g15156(1) = NOR(g13782, g7050)
g22859(1) = AND(g9456, g20734)
g19571(1) = AND(g3498, g16812)
g22172(1) = AND(g8064, g19857)
g15102(1) = NOR(g14591, g6954)
g15127(1) = NOR(g12879, g13605)
g17151(1) = AND(g8659, g12996)
g19752(1) = AND(g2771, g15864)
g15096(1) = NOR(g13191, g12867)
g15116(1) = AND(g4297, g14454)
g21605(1) = AND(g13005, g15695)
g15152(1) = NOR(g13745, g12896)
g16069(2) = NAND(I17447, I17448)
g16893(2) = NAND(g10685, g13252, g703)
g15055(1) = NOR(g6808, g13350)
g15093(1) = NOR(g13177, g6904)
g15164(1) = NOR(g13835, g12906)
g17181(1) = AND(g1945, g13014)
g15130(1) = NOR(g13638, g6985)
g19266(1) = AND(g246, g16214)
g19588(1) = AND(g3849, g16853)
g17699(1) = NAND(I18681, I18682)
g15073(1) = NOR(g12844, g13416)
g19749(1) = AND(g732, g16646)
g22226(1) = OR(g21333, g17655)
g15094(1) = NOR(g13177, g12865)
g15832(1) = NAND(g7903, g7479, g13256)
g19693(1) = AND(g6181, g17087)
g15090(1) = NOR(g13144, g12862)
g15147(1) = NOR(g13716, g12892)
g15109(1) = AND(g4269, g14454)
g20784(1) = NAND(g14616, g17595)
g15108(1) = AND(g4264, g14454)
g15148(1) = NOR(g13716, g12893)
g19914(1) = AND(g2815, g15853)
g17150(1) = AND(g8579, g12995)
g15059(1) = NOR(g12839, g13350)
g15157(1) = NOR(g13782, g12900)
g22217(1) = OR(g21302, g17617)
g19594(1) = AND(g11913, g17268)
g21288(1) = NAND(g14616, g17492)
g17618(1) = NAND(I18580, I18581)
g19637(1) = AND(g5142, g16958)
g15068(1) = NOR(g6826, g13416)
g23151(1) = AND(g18994, g7162)
g21394(1) = AND(g13335, g15799)
g19139(1) = AND(g452, g16195)
g19333(1) = AND(g464, g16223)
g20027(1) = NOR(g16242, g13779)
g20171(1) = AND(g16479, g10476)
g15053(1) = NOR(g12836, g13350)
g19585(1) = AND(g17180, g14004)
g15120(1) = NOR(g12873, g13605)
g15128(1) = NOR(g13638, g12880)
g19674(1) = AND(g2819, g15867)
g19692(1) = AND(g12066, g17086)
g16662(1) = AND(g4552, g14753)
g15113(1) = AND(g4291, g14454)
g15146(1) = NOR(g13716, g7003)
g23103(1) = AND(g10143, g20765)
g15105(1) = AND(g4235, g14454)
g19949(1) = OR(g17671, g14681)
g18893(1) = AND(g16215, g16030)
g15167(1) = NOR(g13835, g12908)
g15088(1) = NOR(g13144, g6874)
g20169(1) = OR(g16184, g13460)
g17179(1) = AND(g1041, g13211)
g15081(1) = AND(g2689, g12983)
g19206(1) = AND(g460, g16206)
g22993(1) = NOR(g1322, g16292, g19873)
g21186(1) = NAND(g14616, g17363)
g15072(1) = NOR(g13416, g12843)
g22762(1) = AND(g9305, g20645)
g20188(1) = AND(g5849, g17772)
g15061(1) = NOR(g6815, g13394)
g19500(1) = AND(g504, g16712)
g20218(1) = AND(g6541, g17815)
g15086(1) = NOR(g13144, g12859)
g15104(1) = AND(g6955, g14454)
g15056(1) = NOR(g6809, g13350)
g21067(1) = AND(g10085, g17625)
g16713(2) = NAND(I17924, I17925)
g23801(1) = AND(g1448, g19362)
g23917(1) = AND(g1472, g19428)
g22720(1) = AND(g9253, g20619)
g22340(1) = AND(g19605, g13522)
g15112(1) = AND(g4284, g14454)
g15097(1) = NOR(g12868, g13191)
g21066(1) = AND(g10043, g17625)
g15141(1) = NOR(g12888, g13680)
g19880(1) = NOR(g16201, g13634)
g23854(1) = AND(g4093, g19506)
g17656(1) = NAND(I18626, I18627)
g17193(1) = AND(g2504, g13023)
g17593(1) = NAND(I18537, I18538)
g18879(1) = OR(g17365, g14423)
g19907(1) = NOR(g16210, g13676)
g15149(1) = NOR(g13745, g12894)
g19906(1) = NOR(g16209, g13672)
g15139(1) = NOR(g12886, g13680)
g19767(1) = AND(g16810, g14203)
g21557(1) = AND(g12980, g15674)
g23405(1) = OR(g19791, g16245)
g17568(1) = NAND(I18486, I18487)
g18906(1) = AND(g13568, g16264)
g19521(1) = AND(g513, g16739)
g15071(1) = NOR(g6831, g13416)
g15080(1) = AND(g12855, g12983)
g20215(1) = AND(g16479, g10476)
g15650(1) = AND(g8362, g13413)
g19462(3) = AND(g7850, g14182, g14177, g16646)
g15087(1) = NOR(g12860, g13144)
g19535(1) = OR(g15651, g13020)
g17091(1) = AND(g8659, g12940)
g23208(1) = NOR(g20035, g16324)
g18934(1) = AND(g3133, g16096)
g17192(1) = AND(g1677, g13022)
g20082(1) = OR(g16026, g13321)
g19661(1) = AND(g5489, g16969)
g19715(1) = AND(g9679, g17120)
g16155(2) = NAND(I17495, I17496)
g22846(1) = AND(g9386, g20676)
g15163(1) = NOR(g13809, g12905)
g17152(1) = AND(g8635, g12997)
g19784(1) = AND(g2775, g15877)
g19354(1) = AND(g471, g16235)
g19575(1) = OR(g15693, g13042)
g18951(1) = AND(g3484, g16124)
g19358(1) = NAND(g15723, g1399)
g19855(1) = AND(g2787, g15962)
g15075(1) = AND(g12850, g12955)
g22304(1) = OR(g21347, g17693)
g15843(1) = NAND(g7922, g7503, g13264)
g16181(1) = NAND(g13475, g13495, g13057, g13459)
g17182(1) = AND(g8579, g13016)
g19384(1) = AND(g667, g16310)
g17624(1) = NAND(I18588, I18589)
g22717(1) = AND(g9291, g20212)
g19735(1) = AND(g9740, g17135)
g15119(1) = AND(g4249, g14454)
g15118(1) = AND(g4253, g14454)
g15066(1) = NOR(g12841, g13394)
g15959(2) = NAND(I17405, I17406)
g21303(1) = AND(g10120, g17625)
g15153(1) = NOR(g13745, g12897)
g20783(1) = NAND(g14616, g17225)
g18981(1) = AND(g11206, g16158)
g19593(1) = OR(g17145, g14210)
g23381(1) = AND(g7239, g21413)
g15150(1) = NOR(g12895, g13745)
g15099(1) = NOR(g13191, g12869)
g15154(1) = NOR(g13782, g12898)
g19660(1) = AND(g12001, g16968)
g11154(1) = NAND(I14212, I14213)
g19655(1) = AND(g2729, g16966)
g15159(1) = NOR(g13809, g12902)
g15095(1) = NOR(g13177, g12866)
g19999(1) = NOR(g16232, g13742)
g19997(1) = NOR(g16231, g13739)
g19487(1) = AND(g499, g16680)
g18950(1) = AND(g11193, g16123)
g15058(1) = NOR(g12838, g13350)
g20051(1) = OR(g15936, g13306)
g19601(1) = AND(g16198, g11149)
g19441(1) = OR(g15507, g12931)
g21405(1) = AND(g13377, g15811)
g21334(1) = NAND(g14616, g17596)
g21187(1) = NAND(g14616, g17364)
g15091(1) = NOR(g13177, g12863)
g15115(1) = AND(g2946, g14454)
g21287(1) = NAND(g14616, g17571)
g19556(1) = AND(g11932, g16809)
g15142(1) = NOR(g13680, g12889)
g15100(1) = NOR(g13191, g12870)
g17199(1) = AND(g2236, g13034)
g22843(1) = AND(g9429, g20272)
g15131(1) = NOR(g12881, g13638)
g19740(1) = AND(g2783, g15907)
g20203(1) = AND(g6195, g17789)
g15064(1) = NOR(g6820, g13394)
g23779(1) = AND(g1105, g19355)
g15155(1) = NOR(g12899, g13782)
g16196(1) = NAND(g13496, g13513, g13079, g13476)
g20063(1) = OR(g15978, g13313)
g15062(1) = NOR(g6817, g13394)
g15051(1) = NOR(g6801, g13350)
g19578(1) = AND(g16183, g11130)
g15132(1) = NOR(g12882, g13638)
g15054(1) = NOR(g12837, g13350)
g15092(1) = NOR(g12864, g13177)
g18987(1) = AND(g182, g16162)
g15114(1) = AND(g4239, g14454)
g15121(1) = NOR(g12874, g13605)
g15082(1) = AND(g2697, g12983)
g15107(1) = AND(g4258, g14454)
g18943(1) = AND(g269, g16099)
g23811(1) = AND(g4087, g19364)
g15098(1) = NOR(g13191, g6927)
g19746(1) = AND(g9816, g17147)
g23412(1) = AND(g7297, g21510)
g19684(1) = AND(g2735, g17297)
g23229(1) = AND(g18994, g4521)
g22309(1) = AND(g1478, g19751)
g22308(1) = AND(g1135, g19738)
g15134(1) = NOR(g13638, g12884)
g18910(1) = AND(g16227, g16075)
g15165(1) = NOR(g12907, g13835)
g15143(1) = NOR(g6998, g13680)
g20034(1) = OR(g15902, g13299)
g22225(1) = OR(g21332, g17654)
g15160(1) = NOR(g12903, g13809)
g19372(1) = AND(g686, g16289)
g15129(1) = NOR(g6984, g13638)
g19335(1) = NAND(g15717, g1056)
g15057(1) = NOR(g6810, g13350)
g19953(1) = NOR(g16220, g13712)
g19951(1) = NOR(g16219, g13709)
g22160(1) = AND(g8005, g19795)
g15123(1) = NOR(g6975, g13605)
g20199(1) = NAND(g16815, g13968, g16749, g13907)
g21363(1) = NAND(g17708, g14664, g17640, g14598)
g20185(1) = NAND(g16772, g13928, g16723, g13882)
g21416(1) = NAND(g17775, g14781, g17744, g14706)
g20134(1) = NAND(g17572, g14542, g17495, g14452)
g20170(1) = NAND(g16741, g13897, g16687, g13866)
g22669(1) = OR(g7763, g19525)
g21357(1) = NAND(g15736, g13109, g15726, g13086)
g21385(1) = NAND(g17736, g14696, g17679, g14636)
g21402(1) = NAND(g17757, g14740, g17716, g14674)
g21365(1) = NAND(g15744, g13119, g15730, g13100)
g20151(1) = NAND(g17598, g14570, g17514, g14519)
g21351(1) = NAND(g15729, g13098, g15720, g13069)
g21433(1) = NAND(g17792, g14830, g17765, g14750)
g21307(1) = NAND(g15719, g13067, g15709, g13040)
g20111(1) = NAND(g17513, g14517, g17468, g14422)
g21339(1) = NAND(g15725, g13084, g15713, g13050)
g16719(1) = NAND(g3243, g13700, g3310, g11350)
g14820(1) = NAND(g6307, g12173, g6315, g12423)
g17761(1) = NAND(g6291, g14529, g6358, g12423)
g14780(1) = NAND(g6275, g12101, g6329, g12423)
g23132(2) = NAND(g8155, g19932)
g23623(2) = NAND(g9364, g20717)
g14686(1) = NAND(g5268, g12059, g5276, g12239)
g16776(1) = NAND(g3945, g13772, g4012, g11419)
g13257(1) = NAND(g1389, g10544)
g17712(1) = NAND(g5599, g14425, g5666, g12301)
g17675(1) = NAND(g5252, g14399, g5320, g12239)
I20487(1) = NAND(g16696, I20486)
I20488(1) = NAND(g16757, I20486)
g23167(2) = NAND(g8219, g19981)
g22306(1) = NAND(g4584, g4616, g13202, g19071)
g13993(1) = NAND(g3961, g11255, g3969, g11419)
g13210(1) = NAND(g7479, g10521)
g13580(2) = NAND(g11849, g7503, g7922, g10544)
g14730(1) = NAND(g5615, g12093, g5623, g12301)
g14695(1) = NAND(g5583, g12029, g5637, g12301)
g14771(1) = NAND(g5961, g12129, g5969, g12351)
g17740(1) = NAND(g5945, g14497, g6012, g12351)
g14739(1) = NAND(g5929, g12067, g5983, g12351)
g23659(2) = NAND(g9434, g20854)
g22709(1) = NAND(g1193, g19611)
g23692(2) = NAND(g9501, g20995)
g11292(2) = NAND(I14331, I14332)
g14829(1) = NAND(g6621, g12137, g6675, g12471)
g22753(1) = NAND(g1536, g19632)
g23079(2) = NOR(g8390, g19965)
I20460(2) = NAND(g17515, g14187)
g21284(2) = NOR(g16646, g9690)
g12332(2) = NAND(I15167, I15168)
g13573(1) = NAND(g8002, g10544, g7582, g1351)
g13058(1) = NAND(g10544, g1312)
g14871(1) = NAND(g6653, g12211, g6661, g12471)
g23642(2) = NOR(g9733, g21124)
g23124(2) = NOR(g8443, g20011)
g20181(1) = NAND(g13252, g16846)
g17779(1) = NAND(g6637, g14556, g6704, g12471)
g13958(1) = NAND(g3610, g11238, g3618, g11389)
g16745(1) = NAND(g3594, g13730, g3661, g11389)
g13927(1) = NAND(g3578, g11207, g3632, g11389)
g13896(1) = NAND(g3227, g11194, g3281, g11350)
g13043(1) = NAND(g10521, g969)
g13967(1) = NAND(g3929, g11225, g3983, g11419)
g14663(1) = NAND(g5236, g12002, g5290, g12239)
g13918(1) = NAND(g3259, g11217, g3267, g11350)
I20468(1) = NAND(g16663, I20467)
I20469(1) = NAND(g16728, I20467)
g23560(2) = NOR(g9607, g20838)
g13240(1) = NAND(g1046, g10521)
g13544(1) = NAND(g7972, g10521, g7549, g1008)
g23105(2) = NAND(g8097, g19887)
g23726(2) = NAND(g9559, g21140)
g13241(1) = NAND(g7503, g10544)
g23602(2) = NOR(g9672, g20979)
g23756(2) = NAND(g9621, g21206)
g23678(2) = NOR(g9809, g21190)
g23711(2) = NOR(g9892, g21253)
g23052(2) = NOR(g8334, g19916)
g13551(2) = NAND(g11812, g7479, g7903, g10521)
g23051(1) = NOR(g7960, g19427)
g23024(1) = NOR(g7936, g19407)
g16349(72) = NOT(I17661)
I19778(1) = NOT(g17781)
g17433(30) = NOT(I18382)
g17821(22) = NOT(I18829)
g17844(1) = NOT(I18832)
g15737(1) = NAND(g13240, g13115, g7903, g13210)
g15426(52) = NOT(I17121)
g17929(22) = NOT(I18855)
g17782(1) = NOT(I18788)
g17062(22) = NOT(I18154)
g17873(52) = NOT(I18849)
g16861(4) = NOT(I18051)
g15348(22) = NOT(I17111)
g15938(20) = NOT(I17401)
g17155(1) = NOT(I18205)
g15563(2) = NOT(I17140)
g18008(52) = NOT(I18868)
g17614(1) = NOT(I18571)
g16777(4) = NOT(I18003)
g18930(1) = NOT(g15789)
g22342(14) = AND(g9354, g9285, g21287)
g16326(22) = NOT(I17658)
g17328(34) = NOT(I18313)
g15748(1) = NAND(g13257, g13130, g7922, g13241)
I20830(1) = NOT(g17657)
g25090(1) = NOT(g23630)
g17428(1) = NOT(I18367)
g24655(1) = NOT(g23067)
g17533(34) = NOT(I18482)
g15573(1) = NOT(I17154)
g15615(12) = NOT(I17181)
g23436(2) = AND(g676, g20375)
g22384(14) = AND(g9354, g9285, g20784)
g15224(52) = NOT(I17101)
g24667(1) = NOT(g23112)
g15277(66) = NOT(I17104)
g16782(12) = NOT(I18006)
g21657(1) = NOT(g17657)
g15373(52) = NOT(I17118)
g16897(22) = NOT(I18083)
g15758(20) = NOT(I17276)
g15171(52) = NOT(I17098)
g17224(1) = NOT(I18248)
I21254(1) = NOT(g16540)
g15509(52) = NOT(I17136)
g16931(22) = NOT(I18101)
g16449(22) = NOT(I17679)
g15634(12) = NOT(I17188)
g17485(1) = NOT(I18408)
g17015(40) = NOT(I18143)
g16508(1) = NOT(I17704)
g16964(1) = NOT(I18120)
g23850(3) = NAND(g12185, g19462)
g25133(1) = NOT(g23733)
g16826(12) = NOT(I18034)
I19857(1) = NOT(g16640)
I18891(1) = NOT(g16676)
g16077(12) = NOT(I17456)
g15595(12) = NOT(I17173)
g21656(1) = NOT(g17700)
g15483(22) = NOT(I17128)
g25255(2) = NAND(g20979, g23659)
g17367(16) = NOT(I18320)
g19592(1) = NOT(I20035)
I21074(1) = NOT(g17766)
I20891(1) = NOT(g17700)
I21238(1) = NOT(g16540)
g17249(14) = NOT(I18265)
g17501(1) = NOT(I18434)
g16971(14) = NOT(I18131)
g16431(16) = NOT(I17675)
g17093(2) = NOT(I18165)
g24685(1) = NOT(g23139)
g16100(18) = NOT(I17471)
I19775(1) = NOT(g17780)
I21722(1) = NOT(g19264)
g23954(1) = NOT(I23099)
g24587(1) = NOT(g23112)
g17096(22) = NOT(I18168)
g17955(52) = NOT(I18865)
I21230(1) = NOT(g16540)
g17125(2) = NOT(I18177)
I20840(1) = NOT(g17727)
I19831(1) = NOT(g16533)
g16987(22) = NOT(I18135)
g16308(1) = NOT(I17636)
g15915(16) = NOT(I17392)
g20230(1) = NOT(I20499)
g17200(12) = NOT(I18238)
g17432(1) = NOT(I18379)
g22417(14) = AND(g7753, g9285, g21186)
g17226(12) = NOT(I18252)
g20060(2) = NOT(g16540)
g21678(2) = NOT(g16540)
g17059(2) = NOT(I18151)
g24579(1) = NOT(g23067)
g16856(4) = NOT(I18048)
g21686(2) = NOT(g16540)
I19843(1) = NOT(g16594)
g15680(12) = NOT(I17207)
g24586(1) = NOT(g23067)
g24842(1) = OR(g7804, g22669)
I18912(1) = NOT(g15050)
g15714(1) = NOT(I17228)
g15569(1) = NOT(I17148)
g17508(1) = NOT(I18443)
I17395(1) = NOT(g12952)
I21013(1) = NOT(g15806)
g16053(12) = NOT(I17442)
g16322(1) = NOT(I17650)
g15656(12) = NOT(I17198)
g20046(2) = NOT(g16540)
g22407(1) = NOT(g19455)
g16923(1) = NOT(I18089)
g17296(1) = NOT(I18280)
g24437(1) = NOT(g22654)
g16136(18) = NOT(I17491)
I19238(1) = NOT(g15079)
g16284(1) = NOT(I17609)
g16877(4) = NOT(I18071)
I20929(1) = NOT(g17663)
g17847(22) = NOT(I18839)
g16489(16) = NOT(I17699)
I20433(1) = NOT(g16234)
I20609(1) = NOT(g16539)
g15979(12) = NOT(I17420)
I20910(1) = NOT(g17197)
I18191(1) = NOT(g14385)
g17327(1) = NOT(I18310)
I19759(1) = NOT(g17767)
I17626(1) = NOT(g14582)
I20569(1) = NOT(g16486)
g20073(2) = NOT(g16540)
I21226(1) = NOT(g16540)
I18245(1) = NOT(g14676)
I20399(1) = NOT(g16205)
g25017(1) = NOT(g23699)
I18897(1) = NOT(g16738)
g17812(1) = NOT(I18810)
g16307(1) = NOT(I17633)
g22457(14) = AND(g7753, g7717, g21288)
g17409(1) = NOT(I18344)
g23620(2) = NOT(I22769)
g24711(1) = NOT(g23139)
g24411(3) = AND(g4584, g22161)
g15345(2) = NOT(I17108)
g15885(16) = NOT(I17374)
g16886(6) = NOT(I18078)
I21234(1) = NOT(g16540)
g22359(1) = NOT(g19495)
g15480(2) = NOT(I17125)
I18304(1) = NOT(g14790)
g18948(1) = NOT(g15800)
g16487(1) = NOT(I17695)
g24814(2) = NAND(g20011, g23167)
g15085(1) = NOT(I17008)
g25016(1) = NOT(g23666)
g16752(4) = NOT(I17976)
g16286(1) = NOT(I17615)
g21653(1) = NOT(g17663)
I20369(1) = NOT(g17690)
g18062(2) = NOT(I18872)
g16601(1) = NOT(I17783)
I17879(1) = NOT(g14386)
g18065(22) = NOT(I18875)
g17271(12) = NOT(I18270)
I20412(1) = NOT(g16213)
g25188(1) = NOT(g23909)
g17326(1) = NOT(I18307)
g22649(1) = NOT(g19063)
g16249(8) = NOT(I17590)
g19869(2) = NOT(g16540)
g25218(1) = NOT(g23949)
I21029(1) = NOT(g15816)
g21674(2) = NOT(g16540)
g22719(1) = NOT(I22024)
I20793(1) = NOT(g17694)
g16031(12) = NOT(I17436)
g15169(1) = NOT(I17094)
I19863(1) = NOT(g16675)
g15733(1) = NOT(I17249)
g17384(4) = NOT(I18323)
g16577(1) = NOT(I17747)
g22472(14) = AND(g7753, g9285, g21289)
I19704(1) = NOT(g17653)
g22498(14) = AND(g7753, g7717, g21334)
g17247(1) = NOT(I18259)
g17926(2) = NOT(I18852)
g17324(1) = NOT(I18301)
g23009(1) = AND(g20196, g14219)
I17557(1) = NOT(g14510)
g16587(1) = NOT(I17763)
g16000(20) = NOT(I17425)
g16821(4) = NOT(I18031)
g25036(1) = NOT(g23733)
g22325(3) = NAND(g1252, g19140)
g16578(1) = NOT(I17750)
g25233(2) = NAND(g20838, g23623)
g17591(1) = NOT(I18526)
g22432(14) = AND(g9354, g7717, g21187)
g24528(3) = NAND(g4098, g22654)
g16309(1) = NOT(I17639)
I21246(1) = NOT(g16540)
g25239(1) = NOT(g23972)
g19954(2) = NOT(g16540)
g24778(1) = NOT(g23286)
g15579(1) = NOT(I17159)
g24809(2) = NAND(g19965, g23132)
g25092(1) = NOT(g23666)
g24999(1) = NOT(g23626)
I19348(1) = NOT(g15084)
g16129(6) = NOT(I17488)
g16816(4) = NOT(I18028)
g15588(1) = NOT(I17166)
g23234(1) = NOT(g20375)
I21058(1) = NOT(g17747)
I18086(1) = NOT(g13856)
g17427(1) = NOT(I18364)
g23782(3) = NAND(g2741, g21062)
g16600(1) = NOT(I17780)
I19484(1) = NOT(g15122)
g17691(1) = NOT(I18674)
g25334(2) = NAND(g21253, g23756)
g24971(1) = NOT(g23590)
I19799(1) = NOT(g17817)
g17952(1) = NOT(I18858)
g17248(1) = NOT(I18262)
I18894(1) = NOT(g16708)
g19446(2) = NOT(I19917)
g21682(2) = NOT(g16540)
g16620(1) = NOT(I17808)
g24484(1) = AND(g16288, g23208)
g22860(1) = NOT(g20000)
g24603(1) = NOT(g23108)
g22497(1) = NOT(g19513)
I18160(1) = NOT(g14441)
g17413(1) = NOT(I18350)
g16164(6) = NOT(I17507)
I19235(1) = NOT(g15078)
I20495(1) = NOT(g16283)
g22527(1) = NOT(g19546)
g17870(1) = NOT(I18842)
I21250(1) = NOT(g16540)
g24626(1) = NOT(g23139)
g22496(1) = NOT(g19510)
g23573(1) = NOT(g20248)
g17818(1) = NOT(I18822)
I19345(1) = NOT(g15083)
g25448(1) = AND(g11202, g22680)
g17590(1) = NOT(I18523)
I22918(1) = NOT(g21451)
I17569(1) = NOT(g14564)
g17526(1) = NOT(I18469)
g16795(4) = NOT(I18009)
g25293(2) = NAND(g21190, g23726)
g23472(1) = NOT(g21062)
g15862(1) = NOT(I17355)
g23716(2) = OR(g9194, g20905)
g16323(1) = NOT(I17653)
g22660(1) = NOT(g19140)
I19012(1) = NOT(g15060)
I18900(1) = NOT(g16767)
g25273(1) = NOT(g23978)
I19789(1) = NOT(g17793)
g17431(1) = NOT(I18376)
I20355(1) = NOT(g17613)
I18414(1) = NOT(g14359)
I21222(1) = NOT(g18091)
g17408(1) = NOT(I18341)
I21042(1) = NOT(g15824)
I18906(1) = NOT(g16963)
g17486(1) = NOT(I18411)
g24985(1) = NOT(g23586)
g19882(2) = NOT(g16540)
I18138(1) = NOT(g14277)
g21659(1) = NOT(g17727)
g17531(1) = NOT(I18476)
g17178(1) = NOT(I18214)
g17953(1) = NOT(I18861)
I18885(1) = NOT(g16643)
g19908(2) = NOT(g16540)
g22369(14) = AND(g9354, g7717, g20783)
I20447(1) = NOT(g16244)
g17587(1) = NOT(I18518)
g23496(1) = NOT(g20248)
I20882(1) = NOT(g17619)
g19866(2) = NOT(g16540)
I21242(1) = NOT(g16540)
g16429(1) = NOT(I17671)
g16428(1) = NOT(I17668)
g17615(1) = NOT(I18574)
I18882(1) = NOT(g16580)
g17430(1) = NOT(I18373)
I21047(1) = NOT(g17429)
I18909(1) = NOT(g16873)
I18114(1) = NOT(g14509)
g21660(1) = NOT(g17694)
g17475(1) = NOT(I18398)
g23550(1) = NOT(g20248)
g19957(2) = NOT(g16540)
g15506(1) = NOT(I17131)
g24665(1) = NOT(g23067)
g21670(2) = NOT(g16540)
g21694(2) = NOT(g16540)
g17128(4) = NOT(I18180)
I17919(1) = NOT(g14609)
g17532(1) = NOT(I18479)
g22408(1) = NOT(g19483)
g21666(2) = NOT(g16540)
g16967(1) = NOT(I18125)
g21654(1) = NOT(g17619)
g23654(1) = NOT(g20248)
g24585(1) = NOT(g23063)
g23192(1) = NOT(g20248)
g25202(1) = NOT(g23932)
g25055(1) = NOT(g23590)
g25111(1) = NOT(g23699)
g25070(1) = NOT(g23590)
I18903(1) = NOT(g16872)
I19851(1) = NOT(g16615)
g23042(3) = NOR(g16581, g19462, g10685)
g17183(4) = NOT(I18221)
g25001(1) = NOT(g23666)
I23149(1) = NOT(g19061)
g17509(1) = NOT(I18446)
g16954(1) = NOT(I18104)
g23578(2) = NOT(I22725)
g24804(2) = NAND(g19916, g23105)
g24683(1) = NOT(g23112)
g16525(1) = NOT(I17723)
I20388(1) = NOT(g17724)
I19734(1) = NOT(g17725)
I19487(1) = NOT(g15125)
I20385(1) = NOT(g16194)
g25131(1) = NOT(g23699)
g17302(4) = NOT(I18285)
g24605(1) = NOT(g23139)
g24795(1) = NOT(g23342)
g23614(1) = NOT(g20248)
g23530(1) = NOT(g20248)
g25015(1) = NOT(g23662)
g16285(1) = NOT(I17612)
g24789(1) = NOT(g23309)
I18888(1) = NOT(g16644)
g15371(1) = NOT(I17114)
g25000(1) = NOT(g23630)
g15566(1) = NOT(I17143)
g24604(1) = NOT(g23112)
g24953(3) = NOR(g10262, g23978, g12259)
g25035(1) = NOT(g23699)
g23204(3) = NOR(g10685, g19462, g16488)
g17188(1) = NOT(I18224)
g22529(1) = NOT(g19549)
g25268(2) = NAND(g21124, g23692)
g21662(2) = NOT(g16540)
g25034(1) = NOT(g23695)
g25153(1) = NOT(g23733)
g23047(2) = NAND(g482, g20000)
g25327(1) = NOT(g22161)
I21258(1) = NOT(g16540)
g25109(1) = NOT(g23666)
g23331(1) = NOT(g20905)
g25174(1) = NOT(g23890)
g24625(1) = NOT(g23135)
g24987(1) = NOT(g23630)
g22312(3) = NAND(g907, g19063)
g25047(1) = NOT(g23733)
g25072(1) = NOT(g23630)
g21690(2) = NOT(g16540)
g22544(1) = NOT(g19589)
g24986(1) = NOT(g23590)
g25046(1) = NOT(g23729)
g23512(1) = NOT(g20248)
g20234(1) = NOR(g17140, g14207)
g22648(1) = OR(g18987, g15652)
g24550(1) = AND(g3684, g23308)
g22588(1) = AND(g79, g20078)
g22832(1) = OR(g19354, g15722)
g24670(1) = AND(g5138, g23590)
g24930(1) = AND(g4826, g23948)
g19401(1) = NOR(g17193, g14296)
g19948(1) = AND(g17515, g16320)
g22625(1) = OR(g18910, g18933)
g22665(1) = AND(g17174, g20905)
g23919(1) = AND(g4122, g19546)
g24410(1) = AND(g3817, g23139)
g25229(1) = AND(g7636, g22654)
g19400(1) = NOR(g17139, g14206)
g19540(1) = AND(g1124, g15904)
g24556(1) = AND(g4035, g23341)
g20084(1) = AND(g11591, g16609)
g24922(1) = AND(g4831, g23931)
g23023(1) = AND(g650, g20248)
g24423(1) = AND(g4950, g22897)
g23275(1) = OR(g19680, g16160)
g24569(1) = AND(g5115, g23382)
g16236(1) = NAND(g13573, g13554, g13058)
g21558(1) = AND(g15904, g13729)
g24639(1) = AND(g6181, g23699)
g24416(1) = AND(g4939, g22870)
g24014(1) = AND(g7933, g19063)
g24430(1) = OR(g23151, g8234)
g19651(1) = AND(g1111, g16119)
g24465(1) = AND(g3827, g23139)
g22538(1) = AND(g14035, g20248)
g23217(1) = OR(g19588, g16023)
g22318(1) = OR(g21394, g17783)
g21419(1) = AND(g16681, g13595)
g22991(1) = AND(g645, g20248)
g24475(1) = AND(g3831, g23139)
g23296(1) = OR(g19691, g16177)
g23836(1) = AND(g4129, g19495)
g24720(1) = NOR(g1322, g23051, g19793)
g22591(1) = OR(g18893, g18909)
g25037(1) = OR(g23103, g19911)
g24790(1) = AND(g7074, g23681)
g24401(1) = OR(g23811, g21298)
g24422(1) = AND(g4771, g22896)
g23298(1) = OR(g19693, g16179)
g24913(1) = AND(g4821, g23908)
g24436(1) = AND(g3125, g23067)
g24607(1) = AND(g5817, g23666)
g24464(1) = AND(g3480, g23112)
g24409(1) = AND(g3484, g23112)
g24606(1) = AND(g5489, g23630)
g19444(1) = NOR(g17192, g14295)
g24796(1) = AND(g7097, g23714)
g23348(1) = AND(g15570, g21393)
g23262(1) = OR(g19661, g16126)
g24757(1) = AND(g7004, g23563)
g23251(1) = OR(g19637, g16098)
g20390(1) = NOR(g17182, g14257)
g22659(1) = OR(g19062, g15673)
g22634(1) = OR(g18934, g15590)
g24820(1) = AND(g13944, g23978)
g20152(1) = AND(g11545, g16727)
g24731(1) = AND(g6519, g23733)
g25285(1) = AND(g22152, g13061)
g24390(1) = OR(g23779, g21285)
g22708(1) = OR(g19266, g15711)
g24640(1) = AND(g6509, g23733)
g19631(1) = AND(g1484, g16093)
g22901(1) = OR(g19384, g15745)
g24482(1) = AND(g6875, g23055)
g22679(1) = OR(g19145, g15701)
g23183(1) = OR(g19545, g15911)
g19534(1) = OR(g15650, g13019)
g23193(1) = OR(g19556, g15937)
g19610(1) = AND(g1141, g16069)
g22684(1) = OR(g19206, g15703)
g19383(1) = AND(g16893, g13223)
g20149(1) = NOR(g17091, g14185)
g24387(1) = AND(g3457, g22761)
g22640(1) = OR(g18951, g15613)
g23920(1) = AND(g4135, g19549)
g24011(1) = AND(g7939, g19524)
g24582(1) = AND(g5808, g23402)
g20112(1) = AND(g13540, g16661)
g24378(1) = AND(g3106, g22718)
g24730(1) = AND(g6177, g23699)
g19613(1) = AND(g1437, g16713)
g19560(3) = AND(g15832, g1157, g10893)
g21251(1) = AND(g13969, g17470)
g16291(1) = NAND(g13551, g13545)
g22641(1) = OR(g18974, g15631)
g24393(1) = AND(g3808, g22844)
g19596(1) = AND(g1094, g16681)
g21420(1) = AND(g16093, g13596)
g16312(1) = NAND(g13580, g13574)
g20602(1) = AND(g10803, g15580)
g22644(1) = OR(g18981, g15632)
g22307(1) = AND(g20027, g21163)
g23197(1) = OR(g19571, g15966)
g23957(1) = AND(g4138, g19589)
g24545(1) = AND(g3333, g23285)
g20977(1) = AND(g10123, g17301)
g22331(1) = OR(g21405, g17809)
g23209(1) = OR(g19585, g19601)
g19568(1) = AND(g1467, g15959)
g22937(1) = AND(g753, g20540)
g22547(2) = OR(g16855, g20215)
g23615(1) = OR(g20109, g20131)
g24495(1) = AND(g6928, g23127)
g24687(1) = AND(g5827, g23666)
g22636(1) = OR(g18943, g15611)
g22653(1) = OR(g18993, g15654)
g24392(1) = AND(g3115, g23067)
g22685(1) = AND(g11891, g20192)
g24488(1) = AND(g6905, g23082)
g24713(1) = AND(g5831, g23666)
g23855(1) = AND(g4112, g19455)
g22216(1) = AND(g13660, g20000)
g24686(1) = AND(g5485, g23630)
g20183(1) = NOR(g17152, g14222)
g22530(1) = OR(g16751, g20171)
g23087(1) = OR(g19487, g15852)
g24589(1) = AND(g5471, g23630)
g22142(1) = AND(g7957, g19140)
g24588(1) = AND(g5142, g23590)
g19788(1) = AND(g9983, g17216)
g23276(1) = OR(g19681, g16161)
g22193(1) = AND(g19880, g20682)
g23885(1) = AND(g4132, g19513)
g24398(1) = OR(g23801, g21296)
g22863(1) = AND(g9547, g20388)
g25366(1) = AND(g7733, g22406)
g23255(1) = OR(g19655, g16122)
g19671(1) = AND(g1454, g16155)
g24008(1) = AND(g7909, g19502)
g23822(1) = OR(g20218, g16929)
g22209(1) = AND(g19907, g20751)
g22208(1) = AND(g19906, g20739)
g23319(1) = OR(g19717, g16193)
g19453(1) = NOR(g17199, g14316)
g23171(1) = OR(g19536, g15903)
g19388(1) = NOR(g17181, g14256)
g23317(1) = OR(g19715, g16191)
g24501(1) = AND(g14000, g23182)
g23884(1) = AND(g4119, g19510)
g24415(1) = AND(g4760, g22869)
g22652(1) = OR(g18992, g15653)
g24608(1) = AND(g6500, g23425)
g23318(1) = OR(g19716, g16192)
g23720(1) = OR(g20165, g16801)
g22751(1) = OR(g19333, g15716)
g24400(1) = AND(g3466, g23112)
g23297(1) = OR(g19692, g16178)
g24443(1) = OR(g23917, g21378)
g23007(1) = AND(g681, g20248)
g24771(1) = AND(g7028, g23605)
g21465(1) = AND(g16155, g13663)
g24432(1) = OR(g23900, g21361)
g24758(1) = AND(g6523, g23733)
g23130(1) = AND(g728, g20248)
g24940(1) = AND(g5011, g23971)
g24399(1) = AND(g3133, g23067)
g19070(1) = NOR(g16957, g11720)
g20135(1) = AND(g16258, g16695)
g23194(1) = OR(g19564, g19578)
g21453(1) = AND(g16713, g13625)
g24580(1) = OR(g22340, g13096)
g19581(3) = AND(g15843, g1500, g10918)
g21464(1) = AND(g16181, g10872)
g24421(1) = AND(g3835, g23139)
g23292(1) = AND(g19879, g16726)
g22662(1) = OR(g19069, g15679)
g21606(1) = AND(g15959, g13763)
g23795(1) = OR(g20203, g16884)
g24649(1) = AND(g6527, g23733)
g24903(1) = AND(g128, g23889)
g19413(1) = NOR(g17151, g14221)
g24395(1) = AND(g4704, g22845)
g23062(1) = AND(g718, g20248)
g23261(1) = OR(g19660, g16125)
g21452(1) = AND(g16119, g13624)
g22299(1) = AND(g19999, g21024)
g22298(1) = AND(g19997, g21012)
g23358(1) = OR(g19746, g16212)
g20162(1) = AND(g8737, g16750)
g24629(1) = AND(g6163, g23699)
g24451(1) = AND(g3476, g23112)
g20628(1) = AND(g1046, g15789)
g24628(1) = AND(g5835, g23666)
g24785(1) = AND(g7051, g23645)
g24557(1) = OR(g22308, g19207)
g24565(1) = OR(g22309, g19275)
g23750(1) = OR(g20174, g16840)
g23374(1) = OR(g19767, g13514)
g22639(1) = OR(g18950, g15612)
g20083(1) = OR(g2902, g17058)
g22664(1) = OR(g19139, g15694)
g24427(1) = AND(g4961, g22919)
g24403(1) = AND(g4894, g22858)
g24572(1) = AND(g5462, g23393)
g23345(1) = OR(g19735, g16203)
g21513(1) = AND(g16196, g10882)
g19430(1) = NOR(g17150, g14220)
g21404(1) = AND(g16069, g13569)
g20095(1) = AND(g8873, g16632)
g24671(1) = AND(g5481, g23630)
g22158(1) = AND(g13698, g19609)
g23153(1) = OR(g19521, g15876)
g23104(1) = AND(g661, g20248)
g24701(1) = NOR(g979, g23024, g19778)
g23770(1) = OR(g20188, g16868)
g24659(1) = AND(g5134, g23590)
g20658(1) = AND(g1389, g15800)
g22645(1) = OR(g18982, g15633)
g23050(1) = AND(g655, g20248)
g20581(1) = AND(g10801, g15571)
g24581(1) = AND(g5124, g23590)
g24714(1) = AND(g6173, g23699)
g24450(1) = AND(g3129, g23067)
g24590(1) = AND(g6154, g23413)
g20094(1) = AND(g8872, g16631)
g23383(1) = OR(g19756, g16222)
g22939(1) = AND(g9708, g21062)
g19436(1) = NOR(g17176, g14233)
g24402(1) = AND(g4749, g22857)
g22219(1) = AND(g19953, g20887)
g22218(1) = AND(g19951, g20875)
g23856(1) = AND(g4116, g19483)
g23346(1) = OR(g19736, g16204)
g16225(1) = NAND(g13544, g13528, g13043)
g23129(1) = OR(g19500, g15863)
g20214(1) = NAND(g16854, g13993, g16776, g13967)
g21384(1) = NAND(g17734, g14686, g17675, g14663)
g20522(1) = OR(g691, g16893)
g21652(1) = NOR(g17619, g17663)
g20198(1) = NAND(g16813, g13958, g16745, g13927)
g21432(1) = NAND(g17790, g14820, g17761, g14780)
g20184(1) = NAND(g16770, g13918, g16719, g13896)
g21401(1) = NAND(g17755, g14730, g17712, g14695)
g21658(1) = NOR(g17694, g17727)
g21655(1) = NOR(g17657, g17700)
g21415(1) = NAND(g17773, g14771, g17740, g14739)
g21462(1) = NAND(g17816, g14871, g17779, g14829)
g19474(1) = NAND(g11609, g17794)
g21353(1) = NAND(g11467, g17157)
g19450(1) = NAND(g11471, g17794)
g21330(1) = NAND(g11401, g17157)
g20076(2) = NAND(g13795, g16521)
g16246(4) = NOR(g13551, g11169)
g20039(1) = NAND(g11250, g17794)
g16272(4) = NOR(g13580, g11189)
g16628(1) = NAND(g3602, g11207, g3618, g13902)
g17581(1) = NAND(g5607, g12029, g5623, g14669)
g21388(1) = NAND(g11608, g17157)
g15787(1) = NAND(g6283, g14575, g6358, g14745)
g15781(1) = NAND(g6267, g12173, g6329, g14745)
g20216(1) = NAND(I20487, I20488)
g21301(1) = NAND(g11371, g17157)
g17608(1) = NAND(g5953, g12067, g5969, g14701)
g20007(1) = NAND(g11512, g17794)
g21294(1) = NAND(g11324, g17157)
g17732(1) = NAND(g3937, g13824, g4012, g13933)
g16604(1) = NAND(g3251, g11194, g3267, g13877)
g20081(1) = NAND(g11325, g17794)
g15741(1) = NAND(g5244, g14490, g5320, g14631)
g21360(1) = NAND(g11510, g17157)
g17650(1) = NAND(g6299, g12101, g6315, g14745)
g25189(2) = NOR(g6082, g23726)
g16660(1) = NAND(g3953, g11225, g3969, g13933)
g24779(2) = NOR(g3736, g23167)
g15734(1) = NAND(g5228, g12059, g5290, g14631)
g25203(2) = NOR(g6428, g23756)
g19466(1) = NAND(g11562, g17794)
g19886(1) = NAND(g11403, g17794)
g24787(1) = NAND(g3391, g23079)
g21345(1) = NAND(g11429, g17157)
I20461(1) = NAND(g17515, I20460)
g15751(1) = NAND(g5591, g14522, g5666, g14669)
I16778(2) = NAND(g11292, g12332)
g24793(1) = NAND(g3742, g23124)
g21359(1) = NAND(g11509, g17157)
g17668(1) = NAND(g3235, g13765, g3310, g13877)
g17634(1) = NAND(g3219, g11217, g3281, g13877)
g21344(1) = NAND(g11428, g17157)
g25200(1) = NAND(g5742, g23642)
g20092(1) = NAND(g11373, g17794)
g17520(1) = NAND(g5260, g12002, g5276, g14631)
g21354(1) = NAND(g11468, g17157)
g24766(2) = NOR(g3385, g23132)
g23324(6) = NAND(g703, g20181)
g21272(1) = NAND(g11268, g17157)
g24776(1) = NAND(g3040, g23052)
g17706(1) = NAND(g3921, g11255, g3983, g13933)
g17689(1) = NAND(g6645, g12137, g6661, g14786)
g20068(1) = NAND(g11293, g17794)
g21377(1) = NAND(g11560, g17157)
g15780(1) = NAND(g5937, g14549, g6012, g14701)
g25237(1) = NAND(g6434, g23711)
g25186(1) = NAND(g5396, g23602)
g21403(1) = NAND(g11652, g17157)
g19962(1) = NAND(g11470, g17794)
g25216(1) = NAND(g6088, g23678)
g20201(1) = NAND(I20468, I20469)
g25172(1) = NAND(g5052, g23560)
g15742(1) = NAND(g5575, g12093, g5637, g14669)
g25175(2) = NOR(g5736, g23692)
g21417(1) = NAND(g11677, g17157)
I20462(1) = NAND(g14187, I20460)
g20055(1) = NAND(g11269, g17794)
g20107(1) = NAND(g11404, g17794)
g21283(1) = NAND(g11291, g17157)
g15752(1) = NAND(g5921, g12129, g5983, g14701)
g25144(2) = NOR(g5046, g23623)
g21331(1) = NAND(g11402, g17157)
g25160(2) = NOR(g5390, g23659)
g24751(2) = NOR(g3034, g23105)
g19442(1) = NAND(g11431, g17794)
g15798(1) = NAND(g6629, g14602, g6704, g14786)
g15788(1) = NAND(g6613, g12211, g6675, g14786)
g17669(1) = NAND(g3570, g11238, g3632, g13902)
g17705(1) = NAND(g3586, g13799, g3661, g13902)
g19913(1) = NAND(g11430, g17794)
g23955(1) = NOR(g2823, g18890)
g23918(1) = NOR(g2799, g21382)
g22190(1) = NOR(g2827, g18949)
g23686(1) = NOR(g2767, g21066)
g23883(1) = NOR(g2779, g21067)
g23871(1) = NOR(g2811, g21348)
g23763(1) = NOR(g2795, g21276)
g23835(1) = NOR(g2791, g21303)
g18092(1) = NOT(I18882)
g18094(1) = NOT(I18888)
g18095(1) = NOT(I18891)
g18096(1) = NOT(I18894)
g18097(1) = NOT(I18897)
g18098(1) = NOT(I18900)
g18099(1) = NOT(I18903)
g18100(1) = NOT(I18906)
g18101(1) = NOT(I18909)
g21894(1) = OR(g20112, g15107)
g24280(1) = OR(g23292, g15109)
g21895(1) = OR(g20135, g15108)
g21891(1) = OR(g19948, g15103)
g18422(1) = NOT(I19238)
g18527(1) = NOT(I19345)
g18093(1) = NOT(I18885)
g18421(1) = NOT(I19235)
g21900(1) = OR(g20977, g15114)
g21896(1) = OR(g20084, g15110)
g21899(1) = OR(g20162, g15113)
g21898(1) = OR(g20152, g15112)
g18528(1) = NOT(I19348)
g21893(1) = OR(g20094, g18655)
g21901(1) = OR(g21251, g15115)
g21897(1) = OR(g20095, g15111)
g21892(1) = OR(g19788, g15104)
g18274(1) = AND(g1311, g16031)
g19635(1) = NOT(g16349)
g20066(1) = NOT(g17433)
g20231(1) = NOT(g17821)
I19786(1) = NOT(g17844)
g21127(10) = NOR(g18065, g12099)
g21308(17) = NOT(g17485)
I20116(1) = NOT(g15737)
g21056(1) = NOT(g15426)
I21210(1) = NOT(g17526)
g19620(7) = NOT(g17296)
g26869(1) = NOT(g24842)
g20511(1) = NOT(g17929)
g25275(6) = NAND(g22342, g11991)
g19606(2) = NOT(g17614)
g19711(1) = NOT(g17062)
g20660(1) = NOT(g17873)
g21461(1) = NOT(g15348)
g19537(1) = NOT(g15938)
g20916(1) = NOT(g18008)
g19492(1) = NOT(g16349)
g25081(1) = NOT(g22342)
g19750(1) = NOT(g16326)
g19984(11) = NOR(g17096, g8171)
g20857(11) = NOR(g17929, g9380)
I20690(1) = NOT(g15733)
g20054(1) = NOT(g17328)
g19919(10) = NOR(g16987, g11205)
I20130(1) = NOT(g15748)
g20773(1) = NOT(I20830)
g20268(1) = NOT(g18008)
g21225(2) = NOT(g17428)
g20180(1) = NOT(g17533)
g20670(1) = NOT(g15426)
g20993(1) = NOT(g15615)
g24839(1) = NOT(g23436)
g24993(1) = NOT(g22384)
g20667(1) = NOT(g15224)
g21069(1) = NOT(g15277)
g21209(11) = NOR(g15483, g9575)
g18975(1) = NOT(g15938)
g19553(1) = NOT(g16782)
I20781(1) = NOT(g17155)
g21068(1) = NOT(g15277)
g18695(1) = AND(g4737, g16053)
g20502(1) = NOT(g15373)
g20210(1) = NOT(g16897)
g19935(11) = NOR(g17062, g8113)
g20618(1) = NOT(g15277)
g21337(1) = NOT(g15758)
g20443(1) = NOT(g15171)
g19757(2) = NOT(g17224)
g18884(1) = NOT(g15938)
g26183(2) = NOR(g23079, g24766)
g18215(1) = AND(g943, g15979)
g21256(10) = NOR(g15483, g12179)
g21425(1) = NOT(g15509)
g20038(1) = NOT(g17328)
g25097(1) = NOT(g22342)
g19673(1) = NOT(g16931)
g21193(10) = NOR(g15348, g12135)
g19397(1) = NOT(g16449)
g21458(1) = NOT(g15758)
g17221(2) = NOT(I18245)
g20601(1) = NOT(g17433)
g21010(1) = NOT(g15634)
g19634(1) = NOT(g16349)
g19872(1) = NOT(g17015)
I20542(1) = NOT(g16508)
I20913(1) = NOT(g16964)
g24791(1) = NOT(g23850)
g25396(2) = NAND(g22384, g2208, g8259)
g20168(1) = NOT(g17533)
g20666(1) = NOT(g15224)
g19574(1) = NOT(g16826)
g19452(1) = NOT(g16326)
g18953(1) = NOT(g16077)
g19912(1) = NOT(g17328)
g21561(1) = NOT(g15595)
g25309(6) = NAND(g22384, g12021)
g21295(1) = NOT(g17533)
g20556(1) = NOT(g15483)
g20580(1) = NOT(g17328)
g26548(1) = NOT(g25255)
g21336(1) = NOT(g17367)
g19780(1) = NOT(g16449)
g26162(2) = NOR(g23052, g24751)
g20110(1) = NOT(g16897)
g20720(11) = NOR(g17847, g9299)
g20922(1) = NOT(I20891)
g20321(1) = NOT(g17821)
g20179(1) = NOT(g17249)
g20178(1) = NOT(g16971)
g19396(1) = NOT(g16431)
g18918(7) = NOT(I19704)
g19731(1) = NOT(g17093)
g20373(1) = NOT(g17929)
g18908(1) = NOT(g16100)
g22139(2) = NOT(I21722)
I24128(1) = NOT(g23009)
g21370(6) = NOT(g16323)
g16677(2) = NOT(I17879)
g20587(1) = NOT(g15373)
g16300(2) = NOT(I17626)
g19787(1) = NOT(g17096)
g20909(1) = NOT(g17955)
g20543(1) = NOT(g17955)
g21669(1) = NOT(I21230)
g19743(1) = NOT(g17125)
g20569(1) = NOT(g15277)
g20568(1) = NOT(g15509)
g19769(1) = NOT(g16987)
g20242(4) = NOT(g16308)
g21424(1) = NOT(g15426)
g21143(11) = NOR(g15348, g9517)
g20772(1) = NOT(g15171)
g19881(1) = NOT(g15915)
g20639(1) = NOT(g15224)
g20638(1) = NOT(g15224)
g20265(1) = NOT(g17821)
g20204(2) = NOT(g16578)
g19662(3) = NOT(g17432)
g21610(1) = NOT(g15615)
I20562(1) = NOT(g16525)
g21189(1) = NOT(g15634)
g24992(1) = NOT(g22417)
g20510(1) = NOT(g17226)
g23189(1) = NOT(g20060)
g25349(6) = NAND(g22432, g12051)
g19482(1) = NOT(g16349)
g20579(1) = NOT(g17249)
g19710(1) = NOT(g17059)
g18983(1) = NOT(g16077)
g19552(1) = NOT(g16856)
g20578(1) = NOT(g15563)
g21383(1) = NOT(g17367)
g19779(1) = NOT(g16431)
g20586(1) = NOT(g15171)
g21267(1) = NOT(g15680)
g20097(2) = NOT(g17691)
g20442(1) = NOT(g15171)
g20086(1) = NOT(I20355)
g19786(1) = NOT(g17062)
g21681(1) = NOT(I21242)
I21115(1) = NOT(g15714)
g20615(1) = NOT(g15509)
g25435(2) = NAND(g22432, g2342, g8316)
g26645(2) = NOR(g23602, g25160)
g20041(4) = NOT(g15569)
g20275(1) = NOT(g17929)
g19968(10) = NOR(g17062, g11223)
g19998(1) = NOT(g15915)
g19672(1) = NOT(g16931)
g21160(2) = NOT(g17508)
g20841(10) = NOR(g17847, g12027)
g21455(1) = NOT(g15426)
g19961(1) = NOT(g17328)
g19505(1) = NOT(g16349)
g21467(1) = NOT(g15758)
g20130(1) = NOT(g17328)
g20998(11) = NOR(g18065, g9450)
g25439(6) = NAND(g22498, g12122)
g20523(1) = NOT(g17821)
g18952(1) = NOT(g16053)
g21352(1) = NOT(g16322)
g21155(1) = NOT(g15656)
g21418(1) = NOT(g17821)
g20006(1) = NOT(g17328)
g19433(1) = NOT(g15915)
g23170(1) = NOT(g20046)
g19387(1) = NOT(g16431)
I20846(1) = NOT(g16923)
g19343(1) = NOT(g16136)
g20703(1) = NOT(g15373)
I21100(1) = NOT(g16284)
g20600(1) = NOT(g15348)
g19368(1) = NOT(g16326)
g20781(1) = NOT(I20840)
g20372(1) = NOT(g17847)
g19412(1) = NOT(g16489)
g20175(2) = NOT(I20433)
g20014(10) = NOR(g17096, g11244)
g25495(2) = NAND(g12483, g22472)
g20516(5) = NOT(I20609)
g18905(1) = NOT(g16077)
g25300(6) = NAND(g22369, g12018)
g21305(1) = NOT(g15758)
g21053(1) = NOT(g15373)
g21466(1) = NOT(g15509)
g21036(1) = NOT(I20910)
g20209(1) = NOT(g17821)
g21560(1) = NOT(g17873)
g20208(1) = NOT(g17533)
g17141(2) = NOT(I18191)
g19379(3) = NOT(g17327)
g25467(2) = NAND(g12432, g22417)
g19050(10) = NOT(I19759)
g20542(1) = NOT(g17873)
I20584(1) = NOT(g16587)
g19386(1) = NOT(g16431)
g20913(1) = NOT(g15373)
g19603(1) = NOT(g16349)
g19742(1) = NOT(g17096)
g20614(1) = NOT(g15426)
g20436(4) = NOT(I20569)
g21693(1) = NOT(I21254)
g20607(1) = NOT(g17955)
g20320(1) = NOT(g17015)
g20274(1) = NOT(g17847)
g20530(1) = NOT(g15509)
g21665(1) = NOT(I21226)
g19338(4) = NOR(g16031, g1306)
g20593(1) = NOT(g15277)
g19429(1) = NOT(g16489)
g18891(1) = NOT(g16053)
g20565(1) = NOT(g18008)
g19730(1) = NOT(g17062)
g19765(1) = NOT(g16897)
g20641(1) = NOT(g15509)
g21454(1) = NOT(g15373)
g19690(1) = NOT(g16826)
g20153(1) = NOT(g16782)
g19504(1) = NOT(g16349)
g20136(7) = NOT(I20399)
g20635(1) = NOT(g18008)
g17010(2) = NOT(I18138)
g20164(1) = NOT(g16826)
g16709(2) = NOT(I17919)
g19128(10) = NOT(I19778)
g21185(1) = NOT(g15277)
g25023(1) = NOT(g22457)
g19626(2) = NOT(g17409)
g17487(1) = NOT(I18414)
g20575(1) = NOT(g17929)
g24474(1) = NOT(g23620)
g20711(1) = NOT(g15509)
g20327(1) = NOT(g15224)
g26830(1) = NOT(g24411)
g26715(2) = NOR(g23711, g25203)
g20537(1) = NOT(g15345)
g19737(1) = NOT(g17015)
I20529(1) = NOT(g16309)
g20606(1) = NOT(g17955)
g19697(1) = NOT(g16886)
g20381(1) = NOT(g17955)
g25385(2) = NAND(g22369, g1783, g8241)
g20091(1) = NOT(g17328)
g21349(1) = NOT(g15758)
g17325(1) = NOT(I18304)
g26093(1) = NOT(g24814)
g18904(1) = NOT(g16053)
g19445(1) = NOT(g15915)
g21304(1) = NOT(g17367)
g19499(1) = NOT(g16782)
g19498(1) = NOT(g16752)
g26686(2) = NOR(g23678, g25189)
g20663(1) = NOT(g15373)
g21139(1) = NOT(g15634)
g21138(1) = NOT(g15634)
g19432(1) = NOT(g15885)
g20553(1) = NOT(g17929)
g20326(1) = NOT(g18008)
g19753(1) = NOT(g16987)
g20536(1) = NOT(g18065)
g20040(1) = NOT(g17271)
g20702(1) = NOT(g17955)
g20904(1) = NOT(g17433)
g19650(1) = NOT(g16971)
g19529(1) = NOT(g16349)
g20564(1) = NOT(g15373)
g19528(1) = NOT(g16349)
g19696(1) = NOT(g17015)
g19330(2) = NOT(g17326)
g18273(1) = AND(g1287, g16031)
g19365(1) = NOT(g16249)
g20673(1) = NOT(g15277)
g21609(1) = NOT(g18008)
g19960(1) = NOT(g17433)
g21608(1) = NOT(g17955)
g20509(1) = NOT(g15277)
g20508(1) = NOT(g15277)
g20634(1) = NOT(g15373)
g21052(1) = NOT(g15373)
g19709(1) = NOT(g16987)
g21463(1) = NOT(g15588)
g19471(1) = NOT(g16449)
g20213(1) = NOT(g17062)
g21184(1) = NOT(g15509)
g20574(1) = NOT(g17847)
g20452(1) = NOT(g17200)
g20912(1) = NOT(g15171)
g19602(1) = NOT(g16349)
g19657(1) = NOT(g16349)
g19068(1) = NOT(g16031)
g19375(1) = NOT(I19863)
g20072(1) = NOT(g17384)
g19878(1) = NOT(g17271)
g20982(10) = NOR(g17929, g12065)
g20592(1) = NOT(g15277)
g21400(1) = NOT(g17847)
g20780(1) = NOT(g15509)
g18929(1) = NOT(g16100)
g21329(1) = NOT(g16577)
g25155(1) = NOT(g22472)
g25170(1) = NOT(g22498)
I19927(1) = NOT(g17408)
g16216(2) = NOT(I17557)
g18827(1) = NOT(g16000)
g25119(1) = NOT(g22384)
g25118(1) = NOT(g22417)
g20583(1) = NOT(g17873)
g19532(1) = NOT(g16821)
g19783(1) = NOT(g16931)
g21414(1) = NOT(g17929)
g21697(1) = NOT(I21258)
g20113(1) = NOT(g16826)
g21407(1) = NOT(g15171)
g19353(1) = NOT(I19831)
g19144(1) = NOT(g16031)
g25101(1) = NOT(g22384)
g20105(1) = NOT(g17433)
g24357(1) = NOT(g22325)
g20640(1) = NOT(g15426)
g20769(1) = NOT(g17955)
g20768(1) = NOT(g17955)
g26518(1) = NOT(g25233)
g25009(1) = NOT(g22472)
g18945(1) = NOT(g16100)
g25008(1) = NOT(g22432)
g20662(1) = NOT(g15171)
g21399(1) = NOT(g15224)
g25892(1) = NOT(g24528)
g21398(1) = NOT(g18008)
g20710(1) = NOT(g15509)
g21278(1) = NOT(I21013)
g20552(1) = NOT(g17847)
g18932(1) = NOT(g16136)
g19687(1) = NOT(g17096)
g20779(1) = NOT(g15509)
g20778(1) = NOT(g15224)
g18897(1) = NOT(g15509)
g21406(1) = NOT(g17955)
g21049(1) = NOT(g17433)
g20380(1) = NOT(g17955)
g26083(1) = NOT(g24809)
g24875(3) = NOR(g8725, g23850, g11083)
g21048(1) = NOT(g17533)
g25154(1) = NOT(g22457)
g20090(1) = NOT(g17433)
g19489(1) = NOT(g16449)
g20233(1) = NOT(g17873)
g20182(1) = NOT(g16897)
g20651(1) = NOT(g15483)
g20672(1) = NOT(g15277)
g21221(1) = NOT(g15680)
g19559(1) = NOT(g16129)
g19558(1) = NOT(g15938)
g25337(2) = NAND(g22342, g1648, g8187)
g20513(1) = NOT(g18065)
g20449(1) = NOT(g15277)
I21006(1) = NOT(g15579)
g19544(1) = NOT(g16349)
g19865(1) = NOT(g15885)
g20448(1) = NOT(g15509)
g19713(1) = NOT(g16816)
g20505(1) = NOT(g15426)
g21689(1) = NOT(I21250)
g20026(1) = NOT(g17271)
g19679(1) = NOT(g16782)
g26209(2) = NOR(g23124, g24779)
g19678(1) = NOT(g16752)
g25083(1) = NOT(g23782)
g19686(1) = NOT(g17062)
I21189(1) = NOT(g17475)
g20433(1) = NOT(g17929)
g18896(1) = NOT(g16031)
g20387(1) = NOT(g15426)
g21421(1) = NOT(g15171)
g26608(1) = NOT(g25334)
g20104(1) = NOT(g17433)
g19890(11) = NOR(g16987, g8058)
g25139(1) = NOT(g22472)
g25138(1) = NOT(g22472)
I19813(1) = NOT(g17952)
g19376(2) = NOT(g17509)
g21434(24) = NOT(g17248)
g21358(1) = NOT(g16307)
g15932(2) = NOT(I17395)
g18944(1) = NOT(g15938)
g20229(1) = NOT(g17015)
g19617(1) = NOT(g16349)
g19470(1) = NOT(g16000)
g19915(1) = NOT(g16349)
g25389(6) = NAND(g22457, g12082)
I22286(1) = NOT(g19446)
g20716(1) = NOT(g15277)
g21291(1) = NOT(g16620)
g19494(1) = NOT(g16349)
g20582(1) = NOT(g17873)
g20627(1) = NOT(g17433)
g20379(1) = NOT(g17821)
g19352(1) = NOT(g15758)
I25028(1) = NOT(g24484)
g20189(1) = NOT(I20447)
g19638(7) = NOT(g17324)
g20386(1) = NOT(g15224)
g18597(1) = AND(g2975, g16349)
g20603(1) = NOT(g17873)
g20096(1) = NOT(g16782)
g17088(2) = NOT(I18160)
I21181(1) = NOT(g17413)
g20681(1) = NOT(g15483)
g19477(1) = NOT(g16431)
g25514(2) = NAND(g12540, g22498)
g20549(1) = NOT(g15277)
g21604(1) = NOT(g15938)
g20548(1) = NOT(g15426)
g20504(1) = NOT(g18008)
g16228(2) = NOT(I17569)
g19748(1) = NOT(g17015)
g19276(1) = NOT(g17367)
g20129(1) = NOT(g17328)
g18880(1) = NOT(g15656)
g21395(1) = NOT(g17873)
g20057(1) = NOT(g16349)
g20128(1) = NOT(g17533)
g20626(1) = NOT(g15483)
g20323(1) = NOT(g17873)
I22289(1) = NOT(g19446)
g20533(1) = NOT(g17271)
g25100(1) = NOT(g22384)
g20775(1) = NOT(g18008)
g18831(1) = NOT(g15224)
g19733(1) = NOT(g16856)
g23777(1) = NOT(I22918)
g20737(1) = NOT(g15656)
g19630(1) = NOT(g16897)
g20232(1) = NOT(g16931)
g25400(6) = NAND(g22472, g12086)
g18989(1) = NOT(g16000)
g21247(1) = NOT(g15171)
g20697(1) = NOT(g17433)
g18988(1) = NOT(g15979)
I25534(1) = NOT(g25448)
g19476(1) = NOT(g16326)
g20512(1) = NOT(g18062)
g19454(1) = NOT(g16349)
g19570(1) = NOT(g16349)
g19712(1) = NOT(g17096)
g21280(1) = NOT(g16601)
g20277(5) = NOT(g16487)
g18887(1) = NOT(g15373)
g20445(1) = NOT(g15224)
I19772(1) = NOT(g17818)
g20499(1) = NOT(g15483)
g21685(1) = NOT(I21246)
g19567(1) = NOT(g16164)
g21061(1) = NOT(I20929)
g20498(1) = NOT(g15348)
g25082(1) = NOT(g22342)
g20611(1) = NOT(g18008)
g20080(1) = NOT(g17328)
I20895(1) = NOT(g16954)
g19519(1) = NOT(g16795)
g19675(1) = NOT(g16987)
g20432(1) = NOT(g17847)
I21067(1) = NOT(g15573)
g20145(1) = NOT(g17533)
g26605(1) = NOT(g25293)
g20650(1) = NOT(g15348)
g20529(1) = NOT(g15509)
g20528(1) = NOT(g15224)
g20696(1) = NOT(g17533)
g25135(1) = NOT(g22457)
g19577(1) = NOT(g16129)
g19439(1) = NOT(g15885)
g20132(1) = NOT(g16931)
g20869(1) = NOT(g15615)
g24960(1) = NOT(g23716)
g19438(1) = NOT(g16249)
g21355(1) = NOT(g17821)
g18878(1) = NOT(g15426)
g20709(1) = NOT(g15426)
g18886(1) = NOT(g16000)
g20127(1) = NOT(I20388)
g20708(1) = NOT(g15426)
g20087(1) = NOT(g17249)
g19566(1) = NOT(g16136)
g18598(1) = AND(g3003, g16349)
g19653(1) = NOT(g16897)
g25341(6) = NAND(g22417, g12047)
g20657(1) = NOT(g17433)
g20774(1) = NOT(g18008)
g19636(1) = NOT(g16987)
g19415(1) = NOT(g15758)
g21059(1) = NOT(g15509)
g19852(1) = NOT(g17015)
g21058(1) = NOT(g15426)
g16960(2) = NOT(I18114)
g19963(1) = NOT(g16326)
g23203(1) = NOT(g20073)
g20994(1) = NOT(g15615)
g24994(1) = NOT(g22432)
g21281(1) = NOT(g16286)
g18977(1) = NOT(g16100)
g19554(1) = NOT(g16861)
g20919(1) = NOT(g15224)
g19200(5) = NOT(I19789)
I21199(1) = NOT(g17501)
g20010(1) = NOT(g17226)
g20918(1) = NOT(g15224)
g18696(1) = AND(g4741, g16053)
g20545(1) = NOT(g15373)
g20079(1) = NOT(g17328)
g20444(1) = NOT(g15373)
g21290(1) = NOT(I21029)
g21156(3) = NOT(g17247)
g20599(1) = NOT(g18065)
g19745(1) = NOT(g16877)
g20598(1) = NOT(g17929)
g19799(1) = NOT(g17062)
g21427(1) = NOT(g17367)
g19798(1) = NOT(g17200)
g20322(1) = NOT(g17873)
g20159(1) = NOT(g17533)
g25121(1) = NOT(g22432)
g20532(1) = NOT(g15277)
g21661(1) = NOT(I21222)
g20158(1) = NOT(g16971)
g19732(1) = NOT(g17096)
g20100(1) = NOT(I20369)
g20561(1) = NOT(g17873)
g20656(1) = NOT(g17249)
g20680(1) = NOT(g15348)
g20144(1) = NOT(g17533)
g19761(1) = NOT(g17015)
g19268(4) = NOR(g15979, g962)
g21297(1) = NOT(I21042)
g19263(1) = NOT(I19799)
g25134(1) = NOT(g22417)
g20631(1) = NOT(g15171)
g18976(1) = NOT(g16100)
g19539(1) = NOT(g16129)
g19773(2) = NOT(g17615)
g18954(2) = NOT(g17427)
g19538(1) = NOT(g16100)
g21181(1) = NOT(g15426)
I19719(1) = NOT(g17431)
g20571(1) = NOT(g15277)
g21222(2) = NOT(g17430)
g21673(1) = NOT(I21234)
g19771(1) = NOT(g17096)
g21426(1) = NOT(g15277)
g20495(1) = NOT(g17926)
g19683(1) = NOT(g16931)
g18830(1) = NOT(g18008)
g20374(1) = NOT(g18065)
g19414(1) = NOT(g16349)
g20669(1) = NOT(g15426)
g20668(1) = NOT(g15426)
g20195(1) = NOT(g16931)
g20525(1) = NOT(g17955)
g18939(1) = NOT(g16077)
g18727(1) = AND(g4931, g16077)
g19367(1) = NOT(I19851)
g18938(1) = NOT(g16053)
g19435(1) = NOT(g16449)
g20544(1) = NOT(g15171)
g20713(1) = NOT(g15277)
g21060(1) = NOT(g15509)
g23060(1) = NOT(g19908)
g18875(1) = NOT(g15171)
g19744(1) = NOT(g15885)
g19345(4) = NOT(g17591)
g25099(1) = NOT(g22369)
g19399(1) = NOT(g16489)
g20610(1) = NOT(g18008)
g21411(1) = NOT(g15426)
g20705(1) = NOT(I20793)
g25098(1) = NOT(g22369)
g19398(1) = NOT(g16489)
g20679(1) = NOT(g15634)
g20270(1) = NOT(g15277)
g19652(1) = NOT(g16897)
g20383(1) = NOT(g15373)
g20267(1) = NOT(g17955)
g25498(2) = NAND(g22498, g2610, g8418)
g19361(1) = NOT(I19843)
g24439(3) = NOR(g7400, g22312)
g21055(1) = NOT(g15224)
g20219(9) = NOT(I20495)
I20937(1) = NOT(g16967)
g18984(2) = NOT(g17486)
g19947(1) = NOT(g17226)
g20617(1) = NOT(g15277)
g19273(1) = NOT(g16100)
g20915(1) = NOT(I20882)
g23019(1) = NOT(g19866)
g19371(1) = NOT(I19857)
g20494(1) = NOT(g17847)
g20623(1) = NOT(g17929)
g20037(1) = NOT(g17328)
g21457(1) = NOT(g17367)
I24400(1) = NOT(g23954)
g20266(1) = NOT(g17873)
g19421(1) = NOT(g16326)
g20853(1) = NOT(g15595)
g21300(1) = NOT(I21047)
g20167(1) = NOT(g16971)
g20194(1) = NOT(g16897)
g20589(1) = NOT(g15224)
g19541(1) = NOT(g16136)
g19473(1) = NOT(g16349)
g20588(1) = NOT(g18008)
g20524(1) = NOT(g17873)
g19789(1) = NOT(g17015)
g25025(1) = NOT(g22498)
g25473(2) = NAND(g12437, g22432)
g19434(1) = NOT(g16326)
g20616(1) = NOT(g15277)
g18874(1) = NOT(g15938)
I19661(1) = NOT(g17587)
g21511(1) = NOT(g15483)
g20704(1) = NOT(g15373)
g20053(1) = NOT(g17328)
g19682(1) = NOT(g17015)
g25120(1) = NOT(g22432)
g18892(1) = NOT(g15680)
g20036(1) = NOT(g17433)
g20101(1) = NOT(g17533)
g20560(1) = NOT(g17328)
g21456(1) = NOT(g15509)
g20642(1) = NOT(g15277)
g26382(3) = NAND(g577, g24953, g12323)
g19760(1) = NOT(g17015)
g18907(1) = NOT(g15979)
g20064(1) = NOT(g17533)
g23085(1) = NOT(g19957)
g20874(1) = NOT(g15680)
g21054(1) = NOT(g15373)
g20630(1) = NOT(g17955)
g21431(1) = NOT(g18065)
g20166(1) = NOT(g16886)
g20009(1) = NOT(g16349)
g20665(1) = NOT(g15373)
g21269(1) = NOT(g15506)
g26625(2) = NOR(g23560, g25144)
g20008(1) = NOT(g16449)
g21268(1) = NOT(g15680)
g19649(1) = NOT(g17015)
g21180(1) = NOT(g18008)
g20555(1) = NOT(g15480)
g19491(1) = NOT(g16349)
g20570(1) = NOT(g15277)
g20712(1) = NOT(g15509)
g20914(1) = NOT(g15373)
g18883(1) = NOT(g15938)
g19755(1) = NOT(g15915)
g19770(1) = NOT(g17062)
g20239(1) = NOT(g17128)
g20567(1) = NOT(g15426)
g20594(1) = NOT(g15277)
g20238(1) = NOT(g17096)
g19794(1) = NOT(g16489)
g19395(1) = NOT(g16431)
g20382(1) = NOT(g15171)
g25429(2) = NAND(g22417, g1917, g8302)
g21279(1) = NOT(g15680)
g19633(1) = NOT(g16931)
g20154(2) = NOT(I20412)
g19719(1) = NOT(g16897)
g20637(1) = NOT(g15224)
g19718(1) = NOT(g17015)
g21286(1) = NOT(g15509)
g19440(1) = NOT(g15915)
g19861(1) = NOT(g17096)
g19573(1) = NOT(g16877)
g21677(1) = NOT(I21238)
g19389(3) = NOT(g17532)
g20501(1) = NOT(g17955)
g20577(1) = NOT(g15483)
I20951(1) = NOT(g17782)
g25024(1) = NOT(g22472)
g19612(1) = NOT(g16897)
g19777(1) = NOT(g17015)
g21410(1) = NOT(g15224)
g20622(1) = NOT(g15595)
g20566(1) = NOT(g15224)
I19707(1) = NOT(g17590)
g19766(1) = NOT(g16449)
g19417(3) = NOT(g17178)
g25852(3) = AND(g4593, g24411)
g18200(1) = NOT(I19012)
g19360(1) = NOT(g16249)
g20636(1) = NOT(g18008)
I19384(1) = NOT(g15085)
g23084(1) = NOT(g19954)
g20852(1) = NOT(g15595)
g21179(1) = NOT(g15373)
g19629(1) = NOT(g17015)
g19451(1) = NOT(g15938)
g21178(1) = NOT(g17955)
g19472(1) = NOT(g16349)
g24963(1) = NOT(g22342)
g20664(1) = NOT(g15373)
g20576(1) = NOT(g18065)
g20585(1) = NOT(g17955)
I23711(1) = NOT(g23192)
g20554(1) = NOT(g15348)
g19776(1) = NOT(g17015)
g19785(1) = NOT(g16987)
g20609(1) = NOT(g15373)
g19754(1) = NOT(g17062)
g20608(1) = NOT(g15171)
g19950(1) = NOT(g15885)
g19370(1) = NOT(g15915)
g20921(1) = NOT(g15426)
g20052(1) = NOT(g17533)
g21423(1) = NOT(g15224)
g19996(1) = NOT(g17271)
g19394(1) = NOT(g16326)
g20674(1) = NOT(g15277)
g20732(1) = NOT(g15595)
g24732(10) = NOT(g23042)
g21123(1) = NOT(g15615)
g18726(1) = AND(g4927, g16077)
g20329(1) = NOT(g15277)
g20207(1) = NOT(g17015)
g20539(1) = NOT(g15483)
g20005(1) = NOT(g17433)
g19902(1) = NOT(g17200)
g24005(2) = NOT(I23149)
g20538(1) = NOT(g15348)
g18991(1) = NOT(g16136)
g19739(1) = NOT(g16931)
g19698(1) = NOT(g16971)
g25157(1) = NOT(g22498)
g20771(1) = NOT(g15171)
g26054(1) = NOT(g24804)
g20235(1) = NOT(g15277)
g19366(1) = NOT(g15885)
g25492(2) = NAND(g12479, g22457)
g20515(1) = NOT(g15483)
g23041(1) = NOT(g19882)
g21275(1) = NOT(g15426)
g24991(1) = NOT(g22369)
g19481(1) = NOT(g16349)
g21340(2) = NOT(I21074)
g19127(1) = NOT(I19775)
g20441(1) = NOT(g17873)
g20584(1) = NOT(g17873)
g19490(1) = NOT(g16489)
g19385(1) = NOT(g16326)
g19980(1) = NOT(g17226)
g20114(12) = NOT(I20385)
g20435(1) = NOT(g15348)
g21362(1) = NOT(g17873)
g24453(3) = NOR(g7446, g22325)
g25156(1) = NOT(g22498)
g19931(1) = NOT(g17200)
g19520(1) = NOT(g16826)
g18947(1) = NOT(g16136)
g19860(1) = NOT(g17226)
g20500(1) = NOT(g17873)
g19659(1) = NOT(g17062)
g20004(1) = NOT(g17249)
g19658(1) = NOT(g16987)
g25039(1) = NOT(g22498)
g20613(1) = NOT(g15224)
g19422(4) = NOR(g16031, g13141)
g19644(4) = NOT(g17953)
g20273(1) = NOT(g17128)
g20106(1) = NOT(g17328)
g20605(1) = NOT(g17955)
g21422(1) = NOT(g15373)
g16920(2) = NOT(I18086)
g24463(1) = NOT(g23578)
g19402(4) = NOR(g15979, g13133)
g19411(1) = NOT(g16489)
g19527(1) = NOT(g16349)
g18829(1) = NOT(g15171)
g19503(1) = NOT(g16349)
g21607(1) = NOT(g17873)
g20514(1) = NOT(g15348)
g18828(1) = NOT(g17955)
g18946(1) = NOT(g16100)
g21274(1) = NOT(g15373)
g20507(1) = NOT(g15509)
g21346(1) = NOT(g17821)
g19714(1) = NOT(g16821)
g26667(2) = NOR(g23642, g25175)
g19979(1) = NOT(g17226)
g20541(1) = NOT(g17821)
g21409(1) = NOT(g18008)
g19741(1) = NOT(g16987)
g21408(1) = NOT(g15373)
g20325(1) = NOT(g15171)
g19067(1) = NOT(g15979)
g20920(1) = NOT(g15426)
g20535(1) = NOT(g17847)
g20434(1) = NOT(g18065)
I20216(1) = NOT(g15862)
g19695(1) = NOT(g17015)
g19526(1) = NOT(g16349)
g18903(1) = NOT(g15758)
g20506(1) = NOT(g15426)
g26823(1) = AND(g24401, g13106)
g20028(4) = NOT(g15371)
g21381(1) = NOT(g18008)
g19689(1) = NOT(g16795)
g25117(1) = NOT(g22417)
g19688(1) = NOT(g16777)
g18990(1) = NOT(g16136)
g18898(4) = NOT(g15566)
g20649(1) = NOT(g18065)
g20240(1) = NOT(g17847)
g20648(1) = NOT(g15615)
g20903(1) = NOT(g17249)
g25432(2) = NAND(g12374, g22384)
g20604(1) = NOT(g17873)
g18832(1) = NOT(g15634)
g19885(1) = NOT(g17249)
g20770(1) = NOT(g17955)
g20563(1) = NOT(g15171)
g19763(1) = NOT(g16431)
g20767(1) = NOT(g17873)
g26340(1) = NOT(g24953)
g21326(2) = NOT(I21058)
g20633(1) = NOT(g15171)
g21252(1) = NOT(g15656)
g19480(1) = NOT(g16349)
g20191(1) = NOT(g17821)
g25007(1) = NOT(g22457)
I19756(1) = NOT(g17812)
g21183(1) = NOT(g15509)
g21397(1) = NOT(g15171)
g19431(1) = NOT(g16249)
g25116(1) = NOT(g22369)
g20573(1) = NOT(g17384)
g20247(1) = NOT(g17015)
g20389(1) = NOT(g15277)
g20612(1) = NOT(g18008)
g20324(1) = NOT(g17955)
g20701(1) = NOT(g17955)
g20777(1) = NOT(g15224)
g20534(1) = NOT(g17183)
g19670(1) = NOT(g16897)
g19734(1) = NOT(g16861)
g19930(1) = NOT(g17200)
g19694(1) = NOT(g16429)
g18911(4) = NOT(g15169)
g21205(1) = NOT(g15656)
g20766(1) = NOT(g17433)
I19796(1) = NOT(g17870)
g21051(1) = NOT(g15171)
g19618(1) = NOT(g16349)
g19443(1) = NOT(g16449)
g20447(1) = NOT(g15426)
g19469(1) = NOT(g16326)
g25006(1) = NOT(g22417)
g19468(1) = NOT(g15938)
g20629(1) = NOT(g17955)
g20451(1) = NOT(g15277)
g21396(1) = NOT(g17955)
g20911(1) = NOT(g15171)
g19677(1) = NOT(g17096)
g20071(1) = NOT(g16826)
g20591(1) = NOT(g15509)
g20776(1) = NOT(g18008)
g25426(2) = NAND(g12371, g22369)
g20147(1) = NOT(g17328)
g25382(2) = NAND(g12333, g22342)
g19410(1) = NOT(g16449)
g24825(9) = NOT(g23204)
g23020(1) = NOT(g19869)
g19479(1) = NOT(g16449)
g19666(3) = NOT(g17188)
g25137(1) = NOT(g22432)
g19478(1) = NOT(g16000)
g18957(16) = NOT(I19734)
g19580(1) = NOT(g16164)
g20446(1) = NOT(g15224)
g20059(1) = NOT(g17302)
g20025(1) = NOT(g17271)
g20058(1) = NOT(g16782)
g19531(1) = NOT(g16816)
g19676(1) = NOT(g17062)
g19685(1) = NOT(g16987)
g19373(1) = NOT(g16449)
g26575(1) = NOT(g25268)
g19654(1) = NOT(g16931)
g18661(1) = NOT(I19487)
g18895(1) = NOT(g16000)
g19800(1) = NOT(g17096)
g20146(1) = NOT(g17533)
g20738(1) = NOT(g15483)
g20562(1) = NOT(g17955)
g21249(1) = NOT(g15509)
g20699(1) = NOT(g17873)
g24699(1) = NOT(g23047)
g21248(1) = NOT(g15224)
g19762(1) = NOT(g16326)
g19964(1) = NOT(g17200)
g20698(1) = NOT(g17873)
g21204(1) = NOT(g15656)
g25136(1) = NOT(g22457)
g20632(1) = NOT(g15171)
g19543(1) = NOT(g16349)
g18889(1) = NOT(g15509)
g18980(1) = NOT(g16136)
g20661(1) = NOT(g15171)
g21380(1) = NOT(g17955)
g20547(1) = NOT(g15224)
g18888(1) = NOT(g15426)
g19569(1) = NOT(g16349)
g19747(1) = NOT(g17015)
g21182(1) = NOT(g15509)
g20715(1) = NOT(g15277)
g20551(1) = NOT(g17302)
g18931(1) = NOT(g16031)
g19772(1) = NOT(g17183)
g20385(1) = NOT(g18008)
g19416(1) = NOT(g15885)
g20103(1) = NOT(g17433)
g24980(1) = NOT(g22384)
g20671(1) = NOT(g15509)
g19579(1) = NOT(g16000)
g19586(1) = NOT(g16349)
g20190(1) = NOT(g16971)
g21343(1) = NOT(g16428)
g25317(3) = NOR(g9766, g23782)
g20546(1) = NOT(g18008)
g20089(1) = NOT(g17533)
g20211(1) = NOT(g16931)
g21369(1) = NOT(g16285)
g20088(1) = NOT(g17533)
g19493(1) = NOT(g16349)
g20497(1) = NOT(g18065)
g21412(1) = NOT(g15758)
g20700(1) = NOT(g17873)
g20659(1) = NOT(g17873)
g20625(1) = NOT(g15348)
g25564(1) = NOT(g22312)
g18894(1) = NOT(g16000)
g21228(24) = NOT(g17531)
g19517(1) = NOT(g16777)
g18979(1) = NOT(g16136)
g19523(1) = NOT(g16100)
g20197(1) = NOT(g16987)
g21379(1) = NOT(g17873)
g18978(1) = NOT(g16000)
g21050(1) = NOT(g17873)
g20527(1) = NOT(g18008)
g25470(2) = NAND(g22457, g2051, g8365)
g19437(1) = NOT(g16349)
g20503(1) = NOT(g15373)
g18877(1) = NOT(g15224)
g18216(1) = AND(g967, g15979)
g20714(1) = NOT(g15277)
g20450(1) = NOT(g15277)
g20707(1) = NOT(g18008)
g21428(1) = NOT(g15758)
g20910(1) = NOT(g15171)
g19600(1) = NOT(g16164)
g19781(1) = NOT(g16489)
g20496(1) = NOT(g17929)
g24979(1) = NOT(g22369)
g19952(1) = NOT(g15915)
g19351(1) = NOT(g17367)
g20978(1) = NOT(g15595)
g24978(1) = NOT(g22342)
g20590(1) = NOT(g15426)
g18917(1) = NOT(g16077)
g19790(1) = NOT(g16971)
g20384(1) = NOT(g18008)
g20067(1) = NOT(g17328)
g25476(2) = NAND(g22472, g2476, g8373)
g21057(1) = NOT(g15426)
g19208(1) = NOT(g17367)
g21299(1) = NOT(g16600)
g20526(1) = NOT(g15171)
g19542(1) = NOT(g16349)
g18102(1) = NOT(I18912)
g20917(1) = NOT(g15224)
g19905(1) = NOT(g15885)
g18876(1) = NOT(g15373)
g18885(1) = NOT(g15979)
g25932(2) = NOR(g7680, g24528)
g19565(1) = NOT(g16000)
g20706(1) = NOT(g18008)
g20597(1) = NOT(g17847)
g20923(1) = NOT(g15277)
g18660(1) = NOT(I19484)
g20624(1) = NOT(g18065)
g19409(1) = NOT(g16431)
g20102(1) = NOT(g17533)
g20157(1) = NOT(g16886)
g18916(1) = NOT(g16053)
g18550(1) = AND(g2819, g15277)
g18314(1) = AND(g1585, g16931)
g18287(1) = AND(g1442, g16449)
g23498(1) = AND(g20234, g12998)
g18307(1) = AND(g1559, g16931)
g18721(1) = AND(g15138, g16077)
g25881(1) = AND(g3821, g24685)
g18596(1) = AND(g2941, g16349)
g18243(1) = AND(g1189, g16431)
g18431(1) = AND(g2185, g18008)
g24763(1) = AND(g17569, g22457)
g18269(1) = AND(g15069, g16031)
g18773(1) = AND(g5694, g15615)
g18341(1) = AND(g1648, g17873)
g18268(1) = AND(g1280, g16000)
g18156(1) = AND(g572, g17533)
g18180(1) = AND(g767, g17328)
g18670(1) = AND(g4621, g15758)
g18734(1) = AND(g4966, g16826)
g18335(1) = AND(g1687, g17873)
g18667(1) = AND(g4601, g17367)
g18694(1) = AND(g4722, g16053)
g18131(1) = AND(g482, g16971)
g24721(1) = AND(g17488, g22369)
g18487(1) = AND(g2441, g15426)
g18619(1) = AND(g3466, g17062)
g18502(1) = AND(g2567, g15509)
g18557(1) = AND(g2771, g15277)
g18210(1) = AND(g936, g15938)
g18618(1) = AND(g3457, g17062)
g18443(1) = AND(g2265, g18008)
g18279(1) = AND(g1361, g16136)
g24813(1) = OR(g22685, g19594)
g18278(1) = AND(g1345, g16136)
g26097(1) = AND(g5821, g25092)
g18469(1) = AND(g2399, g15224)
g18286(1) = AND(g1404, g16164)
g18468(1) = AND(g2393, g15224)
g18306(1) = AND(g15074, g16931)
g25449(1) = AND(g6946, g22496)
g18815(1) = AND(g6523, g15483)
g18601(1) = AND(g3106, g16987)
g18187(1) = AND(g794, g17328)
g18677(1) = AND(g4639, g15758)
g23657(1) = AND(g19401, g11941)
g18143(1) = AND(g586, g17533)
g23428(1) = NAND(g13945, g20522)
g18169(1) = AND(g676, g17433)
g18791(1) = AND(g6044, g15634)
g18168(1) = AND(g681, g17433)
g18410(1) = AND(g2079, g15373)
g18479(1) = AND(g2449, g15426)
g18666(1) = AND(g4593, g17367)
g18363(1) = AND(g1840, g17955)
g18217(1) = AND(g15063, g16100)
g18478(1) = AND(g2445, g15426)
g18486(1) = AND(g2485, g15426)
g18556(1) = AND(g2823, g15277)
g18580(1) = AND(g2907, g16349)
g26050(1) = AND(g9630, g25047)
g18223(1) = AND(g1030, g16100)
g24143(1) = AND(g17694, g21659)
g25368(1) = AND(g6946, g22408)
g26096(1) = AND(g9733, g25268)
g18110(1) = AND(g441, g17015)
g18321(1) = AND(g1620, g17873)
g18179(1) = AND(g763, g17328)
g18531(1) = AND(g2719, g15277)
g18178(1) = AND(g758, g17328)
g18740(1) = AND(g4572, g17384)
g23532(1) = AND(g19400, g11852)
g18186(1) = AND(g753, g17328)
g18676(1) = AND(g4358, g15758)
g18685(1) = AND(g4688, g15885)
g18373(1) = AND(g1890, g15171)
g24015(1) = AND(g19540, g10951)
g18654(1) = AND(g4146, g16249)
g18800(1) = AND(g6187, g15348)
g18417(1) = AND(g2116, g15373)
g18334(1) = AND(g1696, g17873)
g25945(1) = OR(g24427, g22307)
g24990(1) = NOR(g8898, g23324)
g18762(1) = AND(g5475, g17929)
g25050(1) = AND(g13056, g22312)
g18423(1) = AND(g12851, g18008)
g18587(1) = AND(g2980, g16349)
g18543(1) = AND(g2779, g15277)
g26323(1) = AND(g10262, g25273)
g24676(1) = AND(g2748, g23782)
g18117(1) = AND(g464, g17015)
g25802(1) = AND(g8106, g24586)
g18569(1) = AND(g94, g16349)
g18568(1) = AND(g37, g16349)
g18747(1) = AND(g5138, g17847)
g18242(1) = AND(g962, g16431)
g18123(1) = AND(g479, g16886)
g18814(1) = AND(g6519, g15483)
g24762(1) = AND(g655, g23573)
g18751(1) = AND(g5156, g17847)
g18807(1) = AND(g6386, g15656)
g18772(1) = AND(g5689, g15615)
g18639(1) = AND(g3831, g17096)
g18230(1) = AND(g1111, g16326)
g18293(1) = AND(g1484, g16449)
g18638(1) = AND(g3827, g17096)
g18265(1) = AND(g1270, g16000)
g18416(1) = AND(g2112, g15373)
g18391(1) = AND(g1982, g15171)
g18510(1) = AND(g2625, g15509)
g25323(1) = AND(g6888, g22359)
g18579(1) = AND(g2984, g16349)
g24747(1) = AND(g17510, g22417)
g21559(1) = AND(g16236, g10897)
g18578(1) = AND(g2873, g16349)
g18586(1) = AND(g2886, g16349)
g24935(1) = OR(g22937, g19749)
g18442(1) = AND(g2259, g18008)
g25941(1) = OR(g24416, g22219)
g18116(1) = AND(g168, g17015)
g18615(1) = AND(g3347, g17200)
g18720(1) = AND(g15137, g16795)
g25880(1) = AND(g8443, g24814)
g18275(1) = AND(g15070, g16136)
g26145(1) = AND(g11962, g25131)
g18430(1) = AND(g2204, g18008)
g18746(1) = AND(g5134, g17847)
g18493(1) = AND(g2514, g15426)
g18465(1) = AND(g2384, g15224)
g18237(1) = AND(g1146, g16326)
g18340(1) = AND(g1720, g17873)
g18806(1) = AND(g6381, g15656)
g18684(1) = AND(g4681, g15885)
g18142(1) = AND(g577, g17533)
g18517(1) = AND(g2652, g15509)
g25988(1) = AND(g9510, g25016)
g24976(1) = NOR(g671, g23324)
g18130(1) = AND(g528, g16971)
g18193(1) = AND(g837, g17821)
g18362(1) = AND(g1834, g17955)
g20200(1) = NAND(I20461, I20462)
g18165(1) = AND(g650, g17433)
g18523(1) = AND(g2675, g15509)
g26087(1) = AND(g5475, g25072)
g18475(1) = AND(g12853, g15426)
g18222(1) = AND(g1024, g16100)
g18437(1) = AND(g2241, g18008)
g24142(1) = AND(g17700, g21657)
g18703(1) = AND(g4776, g16782)
g18347(1) = AND(g1756, g17955)
g18253(1) = AND(g1211, g16897)
g18600(1) = AND(g3111, g16987)
g18781(1) = AND(g5831, g18065)
g18236(1) = AND(g15065, g16326)
g18351(1) = AND(g1760, g17955)
g18372(1) = AND(g1886, g15171)
g18175(1) = AND(g744, g17328)
g18821(1) = AND(g15168, g15680)
g18264(1) = AND(g1263, g16000)
g18790(1) = AND(g6040, g15634)
g18137(1) = AND(g538, g17249)
g18516(1) = AND(g2638, g15509)
g26078(1) = AND(g5128, g25055)
g24703(1) = AND(g17592, g22369)
g18209(1) = AND(g921, g15938)
g26086(1) = AND(g9672, g25255)
g18208(1) = AND(g930, g15938)
g25879(1) = AND(g11135, g24683)
g18542(1) = AND(g2787, g15277)
g18453(1) = AND(g2315, g15224)
g18614(1) = AND(g3343, g17200)
g18436(1) = AND(g2227, g18008)
g25967(1) = AND(g9373, g24986)
g18607(1) = AND(g3139, g16987)
g18320(1) = AND(g1616, g17873)
g18530(1) = AND(g2715, g15277)
g18593(1) = AND(g2999, g16349)
g18346(1) = AND(g1752, g17955)
g20056(1) = AND(g16291, g9007, g8954, g8903)
g18122(1) = AND(g15052, g17015)
g18565(1) = AND(g2852, g16349)
g18464(1) = AND(g2370, g15224)
g18641(1) = AND(g3841, g17096)
g18797(1) = AND(g6173, g15348)
g18292(1) = AND(g1472, g16449)
g18153(1) = AND(g626, g17533)
g18409(1) = AND(g2084, g15373)
g18136(1) = AND(g550, g17249)
g18408(1) = AND(g2070, g15373)
g18635(1) = AND(g3808, g17096)
g26023(1) = AND(g9528, g25036)
g18164(1) = AND(g699, g17433)
g18575(1) = AND(g2878, g16349)
g18474(1) = AND(g2287, g15224)
g18711(1) = AND(g15136, g15915)
g18327(1) = AND(g1636, g17873)
g22872(1) = OR(g19372, g19383)
g18109(1) = AND(g437, g17015)
g18537(1) = AND(g6856, g15277)
g18108(1) = AND(g433, g17015)
g25966(1) = AND(g9364, g24985)
g18283(1) = AND(g1384, g16136)
g18606(1) = AND(g3133, g16987)
g18492(1) = AND(g2523, g15426)
g18303(1) = AND(g1536, g16489)
g23989(1) = OR(g20581, g17179)
g18750(1) = AND(g15145, g17847)
g18381(1) = AND(g1882, g15171)
g18174(1) = AND(g739, g17328)
g18796(1) = AND(g6167, g15348)
g18390(1) = AND(g1978, g15171)
g18192(1) = AND(g817, g17821)
g25816(1) = AND(g8164, g24604)
g25447(1) = NOR(g23883, g14645)
g18522(1) = AND(g2671, g15509)
g18663(1) = AND(g4311, g17367)
g25976(1) = AND(g9443, g25000)
g23577(1) = AND(g19444, g13033)
g18483(1) = AND(g2453, g15426)
g24750(1) = AND(g17662, g22472)
g18553(1) = AND(g2827, g15277)
g18326(1) = AND(g1664, g17873)
g18536(1) = AND(g2748, g15277)
g18702(1) = AND(g15133, g16856)
g18757(1) = AND(g5352, g15595)
g18252(1) = AND(g990, g16897)
g18621(1) = AND(g3476, g17062)
g25559(1) = AND(g13004, g22649)
g18564(1) = AND(g2844, g16349)
g18183(1) = AND(g781, g17328)
g18673(1) = AND(g4643, g15758)
g18397(1) = AND(g2004, g15373)
g18509(1) = AND(g2587, g15509)
g18508(1) = AND(g2606, g15509)
g18634(1) = AND(g3813, g17096)
g24702(1) = AND(g17464, g22342)
g18213(1) = AND(g952, g15979)
g25938(1) = AND(g8997, g24953)
g18574(1) = AND(g2882, g16349)
g18452(1) = AND(g2311, g15224)
g18205(1) = AND(g904, g15938)
g23554(1) = AND(g20390, g13024)
g18311(1) = AND(g1554, g16931)
g25875(1) = AND(g8390, g24809)
g18592(1) = AND(g2994, g16349)
g18756(1) = AND(g5348, g15595)
g18780(1) = AND(g5827, g18065)
g25929(1) = OR(g24395, g22193)
g18350(1) = AND(g1779, g17955)
g18820(1) = AND(g15166, g15563)
g18152(1) = AND(g613, g17533)
g18396(1) = AND(g2008, g15373)
g18731(1) = AND(g15140, g16861)
g18413(1) = AND(g2089, g15373)
g26119(1) = AND(g11944, g25109)
g18691(1) = AND(g4727, g16053)
g18405(1) = AND(g2040, g15373)
g18583(1) = AND(g2936, g16349)
g25521(1) = NOR(g23955, g14645)
g18113(1) = AND(g405, g17015)
g18787(1) = AND(g15158, g15634)
g18282(1) = AND(g1379, g16136)
g18302(1) = AND(g1514, g16489)
g18357(1) = AND(g1816, g17955)
g18105(1) = AND(g417, g17015)
g18743(1) = AND(g5115, g17847)
g18640(1) = AND(g3835, g17096)
g18769(1) = AND(g15151, g18062)
g18768(1) = AND(g5503, g17929)
g18803(1) = AND(g15161, g15480)
g18662(1) = AND(g15126, g17367)
g18249(1) = AND(g1216, g16897)
g18482(1) = AND(g2472, g15426)
g18248(1) = AND(g15067, g16897)
g18710(1) = AND(g15135, g17302)
g18552(1) = AND(g2815, g15277)
g18204(1) = AND(g914, g15938)
g18779(1) = AND(g5821, g18065)
g18778(1) = AND(g5817, g18065)
g25874(1) = AND(g11118, g24665)
g18786(1) = AND(g15156, g15345)
g18647(1) = AND(g4040, g17271)
g18356(1) = AND(g1802, g17955)
g18826(1) = AND(g7097, g15680)
g18380(1) = AND(g1926, g15171)
g18233(1) = AND(g1094, g16326)
g18182(1) = AND(g776, g17328)
g18651(1) = AND(g15102, g16249)
g18672(1) = AND(g15127, g15758)
g25789(1) = OR(g25285, g14543)
g26089(1) = OR(g24501, g22534)
g18331(1) = AND(g1682, g17873)
g18513(1) = AND(g2575, g15509)
g18449(1) = AND(g12852, g15224)
g18448(1) = AND(g2153, g18008)
g18505(1) = AND(g2583, g15509)
g18404(1) = AND(g2066, g15373)
g24786(1) = AND(g661, g23654)
g18717(1) = AND(g4849, g15915)
g18212(1) = AND(g947, g15979)
g24651(1) = AND(g2741, g23472)
g18723(1) = AND(g4922, g16077)
g18149(1) = AND(g608, g17533)
g18433(1) = AND(g2197, g18008)
g18387(1) = AND(g1955, g15171)
g18620(1) = AND(g3470, g17062)
g18148(1) = AND(g562, g17533)
g18104(1) = AND(g392, g17015)
g18811(1) = AND(g6500, g15483)
g18646(1) = AND(g4031, g17271)
g18343(1) = AND(g12847, g17955)
g18369(1) = AND(g12848, g15171)
g18368(1) = AND(g1728, g17955)
g18412(1) = AND(g2098, g15373)
g18133(1) = AND(g15055, g17249)
g23514(1) = AND(g20149, g11829)
g24723(1) = AND(g17490, g22384)
g18229(1) = AND(g1099, g16326)
g18228(1) = AND(g1061, g16129)
g18716(1) = AND(g4878, g15915)
g18582(1) = AND(g2922, g16349)
g18310(1) = AND(g1333, g16931)
g25247(1) = NOR(g23763, g14645)
g18627(1) = AND(g15093, g17093)
g18379(1) = AND(g1906, g15171)
g18112(1) = AND(g182, g17015)
g18378(1) = AND(g1932, g15171)
g18386(1) = AND(g1964, g15171)
g18603(1) = AND(g3119, g16987)
g18742(1) = AND(g5120, g17847)
g18681(1) = AND(g4653, g15885)
g18802(1) = AND(g6195, g15348)
g18429(1) = AND(g2193, g18008)
g18730(1) = AND(g4950, g16861)
g18793(1) = AND(g6159, g15348)
g18428(1) = AND(g2169, g18008)
g18765(1) = AND(g5489, g17929)
g18690(1) = AND(g15130, g16053)
g18549(1) = AND(g2799, g15277)
g18548(1) = AND(g2807, g15277)
g18504(1) = AND(g2579, g15509)
g18317(1) = AND(g12846, g17873)
g18129(1) = AND(g518, g16971)
g18128(1) = AND(g504, g16971)
g18245(1) = AND(g1193, g16431)
g18626(1) = AND(g3498, g17062)
g18323(1) = AND(g1632, g17873)
g18299(1) = AND(g1526, g16489)
g18533(1) = AND(g2729, g15277)
g24765(1) = AND(g17699, g22498)
g18298(1) = AND(g15073, g16489)
g18775(1) = AND(g7028, g15615)
g18737(1) = AND(g4975, g16826)
g18232(1) = AND(g1124, g16326)
g18697(1) = AND(g4749, g16777)
g18261(1) = AND(g1256, g16000)
g24002(1) = AND(g19613, g10971)
g18512(1) = AND(g2619, g15509)
g23990(1) = AND(g19610, g10951)
g18445(1) = AND(g2273, g18008)
g24775(1) = AND(g17594, g22498)
g18499(1) = AND(g2476, g15426)
g18316(1) = AND(g1564, g16931)
g18498(1) = AND(g2547, g15426)
g18611(1) = AND(g15090, g17200)
g18722(1) = AND(g4917, g16077)
g18432(1) = AND(g2223, g18008)
g18271(1) = AND(g1296, g16031)
g18753(1) = AND(g15148, g15595)
g18461(1) = AND(g2307, g15224)
g18342(1) = AND(g1592, g17873)
g18145(1) = AND(g582, g17533)
g18199(1) = AND(g832, g17821)
g18650(1) = AND(g6928, g17271)
g18736(1) = AND(g4991, g16826)
g18198(1) = AND(g15059, g17821)
g18529(1) = AND(g2712, g15277)
g18330(1) = AND(g1668, g17873)
g18393(1) = AND(g1917, g15171)
g24498(1) = AND(g14036, g23850)
g26049(1) = AND(g9621, g25046)
g18764(1) = AND(g5485, g17929)
g18365(1) = AND(g1848, g17955)
g18132(1) = AND(g513, g16971)
g24722(1) = AND(g17618, g22417)
g18161(1) = AND(g691, g17433)
g18709(1) = AND(g59, g17302)
g18259(1) = AND(g15068, g16000)
g18225(1) = AND(g1041, g16100)
g18708(1) = AND(g4818, g16782)
g25804(1) = AND(g8069, g24587)
g18471(1) = AND(g2407, g15224)
g18258(1) = AND(g1221, g16897)
g18244(1) = AND(g1171, g16431)
g25962(1) = AND(g9258, g24971)
g24764(1) = AND(g17570, g22472)
g18602(1) = AND(g3115, g16987)
g18810(1) = AND(g6505, g15483)
g18657(1) = AND(g4308, g17128)
g18774(1) = AND(g5698, g15615)
g18375(1) = AND(g1902, g15171)
g25833(1) = AND(g8228, g24626)
g18337(1) = AND(g1706, g17873)
g18171(1) = AND(g728, g17433)
g18792(1) = AND(g7051, g15634)
g23996(1) = AND(g19596, g10951)
g18459(1) = AND(g2331, g15224)
g18425(1) = AND(g2161, g18008)
g18458(1) = AND(g2357, g15224)
g20069(1) = AND(g16312, g9051, g9011, g8955)
g18545(1) = AND(g2783, g15277)
g24500(1) = OR(g24011, g21605)
g18444(1) = AND(g2269, g18008)
g24774(1) = AND(g718, g23614)
g18599(1) = AND(g2955, g16349)
g26121(1) = AND(g6167, g25111)
g18817(1) = AND(g6533, g15483)
g18322(1) = AND(g1608, g17873)
g18159(1) = AND(g671, g17433)
g18125(1) = AND(g15053, g16886)
g18532(1) = AND(g2724, g15277)
g18158(1) = AND(g667, g17433)
g18783(1) = AND(g5841, g18065)
g18561(1) = AND(g2841, g15277)
g18656(1) = AND(g15120, g17128)
g18353(1) = AND(g1772, g17955)
g18295(1) = AND(g1489, g16449)
g18680(1) = AND(g15128, g15885)
g18144(1) = AND(g590, g17533)
g18823(1) = AND(g6727, g15680)
g18336(1) = AND(g1700, g17873)
g25936(1) = OR(g24403, g22209)
g25788(1) = AND(g8010, g24579)
g18631(1) = AND(g3694, g17226)
g18364(1) = AND(g1844, g17955)
g24496(1) = OR(g24008, g21557)
g18289(1) = AND(g1448, g16449)
g18309(1) = AND(g1339, g16931)
g18288(1) = AND(g1454, g16449)
g18224(1) = AND(g1036, g16100)
g18571(1) = AND(g2856, g16349)
g18308(1) = AND(g6832, g16931)
g24144(1) = AND(g17727, g21660)
g23551(1) = AND(g10793, g18948)
g18495(1) = AND(g2533, g15426)
g18816(1) = AND(g6527, g15483)
g18687(1) = AND(g4664, g15885)
g22143(1) = AND(g19568, g10971)
g24391(1) = NOR(g22190, g14645)
g18752(1) = AND(g15146, g17926)
g18374(1) = AND(g1878, g15171)
g18643(1) = AND(g3849, g17096)
g18669(1) = AND(g4608, g17367)
g25004(1) = NOR(g676, g23324)
g18260(1) = AND(g1252, g16000)
g18668(1) = AND(g4322, g17367)
g18392(1) = AND(g1988, g15171)
g18195(1) = AND(g847, g17821)
g18489(1) = AND(g2509, g15426)
g18559(1) = AND(g12856, g15277)
g18525(1) = AND(g2610, g15509)
g18488(1) = AND(g2495, g15426)
g18424(1) = AND(g2165, g18008)
g18558(1) = AND(g2803, g15277)
g18544(1) = AND(g2791, g15277)
g18713(1) = AND(g4836, g15915)
g18610(1) = AND(g15088, g17059)
g18705(1) = AND(g4801, g16782)
g25990(1) = AND(g9461, g25017)
g18255(1) = AND(g1087, g16897)
g18189(1) = AND(g812, g17821)
g18679(1) = AND(g4633, g15758)
g18270(1) = AND(g1291, g16031)
g18188(1) = AND(g807, g17328)
g18124(1) = AND(g102, g16886)
g18678(1) = AND(g66, g15758)
g18460(1) = AND(g2351, g15224)
g18686(1) = AND(g4659, g15885)
g18383(1) = AND(g1950, g15171)
g25832(1) = AND(g8219, g24625)
g18267(1) = AND(g1266, g16000)
g18294(1) = AND(g15072, g16449)
g25005(1) = NOR(g6811, g23324)
g18219(1) = AND(g969, g16100)
g25935(1) = OR(g24402, g22208)
g18218(1) = AND(g1008, g16100)
g18160(1) = AND(g645, g17433)
g18455(1) = AND(g2327, g15224)
g18617(1) = AND(g3462, g17062)
g18470(1) = AND(g2403, g15224)
g23581(1) = AND(g20183, g11900)
g18201(1) = AND(g15061, g15938)
g18277(1) = AND(g1312, g16136)
g26147(1) = AND(g6513, g25133)
g25871(1) = AND(g8334, g24804)
g18595(1) = AND(g2927, g16349)
g18467(1) = AND(g2380, g15224)
g18494(1) = AND(g2527, g15426)
g18623(1) = AND(g3484, g17062)
g18782(1) = AND(g5835, g18065)
g25261(1) = OR(g23348, g20193)
g18419(1) = AND(g2051, g15373)
g18352(1) = AND(g1798, g17955)
g18155(1) = AND(g15056, g17533)
g18418(1) = AND(g2122, g15373)
g18822(1) = AND(g6723, g15680)
g18266(1) = AND(g1274, g16000)
g18170(1) = AND(g661, g17433)
g18167(1) = AND(g718, g17433)
g18194(1) = AND(g843, g17821)
g18589(1) = AND(g2902, g16349)
g18588(1) = AND(g2970, g16349)
g18524(1) = AND(g2681, g15509)
g24467(1) = AND(g13761, g23047)
g18401(1) = AND(g2036, g15373)
g18477(1) = AND(g2429, g15426)
g18119(1) = AND(g475, g17015)
g18118(1) = AND(g471, g17015)
g18749(1) = AND(g5148, g17847)
g18616(1) = AND(g6875, g17200)
g18313(1) = AND(g1430, g16931)
g26120(1) = AND(g9809, g25293)
g18748(1) = AND(g5142, g17847)
g25367(1) = AND(g6946, g22407)
g18276(1) = AND(g1351, g16136)
g18285(1) = AND(g1395, g16164)
g26146(1) = AND(g9892, g25334)
g18704(1) = AND(g4793, g16782)
g18305(1) = AND(g1521, g16489)
g18254(1) = AND(g1236, g16897)
g18809(1) = AND(g7074, g15656)
g18466(1) = AND(g2389, g15224)
g18808(1) = AND(g6390, g15656)
g18177(1) = AND(g749, g17328)
g18560(1) = AND(g2837, g15277)
g18642(1) = AND(g15097, g17096)
g18733(1) = AND(g15141, g16877)
g24749(1) = AND(g17511, g22432)
g18630(1) = AND(g3689, g17226)
g18693(1) = AND(g4717, g16053)
g24748(1) = AND(g17656, g22457)
g18166(1) = AND(g655, g17433)
g18665(1) = AND(g4584, g17367)
g24704(1) = AND(g17593, g22384)
g18476(1) = AND(g2433, g15426)
g18485(1) = AND(g2465, g15426)
g18555(1) = AND(g2834, g15277)
g18454(1) = AND(g2303, g15224)
g18570(1) = AND(g2848, g16349)
g18712(1) = AND(g4843, g15915)
g26095(1) = AND(g11923, g25090)
g18239(1) = AND(g1135, g16326)
g18567(1) = AND(g2894, g16349)
g18594(1) = AND(g12858, g16349)
g18238(1) = AND(g1152, g16326)
g24630(1) = AND(g23255, g14149)
g18382(1) = AND(g1936, g15171)
g24009(1) = AND(g19671, g10971)
g18519(1) = AND(g2648, g15509)
g18176(1) = AND(g732, g17328)
g18185(1) = AND(g790, g17328)
g18675(1) = AND(g4349, g15758)
g18518(1) = AND(g2657, g15509)
g18154(1) = AND(g622, g17533)
g18637(1) = AND(g3821, g17096)
g18501(1) = AND(g12854, g15509)
g18729(1) = AND(g15139, g16821)
g18577(1) = AND(g2988, g16349)
g23619(1) = AND(g19453, g13045)
g18728(1) = AND(g4939, g16821)
g18439(1) = AND(g2250, g18008)
g23618(1) = AND(g19388, g11917)
g18438(1) = AND(g2236, g18008)
g24675(1) = AND(g17568, g22342)
g18349(1) = AND(g1768, g17955)
g18348(1) = AND(g1744, g17955)
g18284(1) = AND(g15071, g16164)
g18304(1) = AND(g1542, g16489)
g18622(1) = AND(g3480, g17062)
g18566(1) = AND(g2860, g16349)
g18139(1) = AND(g542, g17249)
g18653(1) = AND(g4176, g16249)
g18138(1) = AND(g546, g17249)
g18636(1) = AND(g3817, g17096)
g18415(1) = AND(g2108, g15373)
g18333(1) = AND(g1691, g17873)
g25987(1) = AND(g9501, g25015)
g18664(1) = AND(g4332, g17367)
g18576(1) = AND(g2868, g16349)
g18585(1) = AND(g2960, g16349)
g18484(1) = AND(g2491, g15426)
g25969(1) = AND(g9310, g24987)
g18554(1) = AND(g2831, g15277)
g18609(1) = AND(g3147, g16987)
g24139(1) = AND(g17619, g21653)
g18312(1) = AND(g1579, g16931)
g18608(1) = AND(g15087, g16987)
g18115(1) = AND(g460, g17015)
g18745(1) = AND(g5128, g17847)
g18799(1) = AND(g6181, g15348)
g23531(1) = AND(g10760, g18930)
g18813(1) = AND(g6513, g15483)
g25503(1) = AND(g6888, g22529)
g18798(1) = AND(g6177, g15348)
g18184(1) = AND(g785, g17328)
g18805(1) = AND(g6377, g15656)
g18674(1) = AND(g4340, g15758)
g25450(1) = AND(g6888, g22497)
g18732(1) = AND(g4961, g16877)
g22490(1) = OR(g21513, g12795)
g25818(1) = AND(g8124, g24605)
g24517(1) = OR(g22158, g18906)
g18692(1) = AND(g4732, g16053)
g18761(1) = AND(g5471, g17929)
g25978(1) = AND(g9391, g25001)
g18400(1) = AND(g2012, g15373)
g26077(1) = AND(g9607, g25233)
g24745(1) = AND(g650, g23550)
g18214(1) = AND(g939, g15979)
g18329(1) = AND(g1612, g17873)
g18207(1) = AND(g925, g15938)
g18539(1) = AND(g2763, g15277)
g18328(1) = AND(g1657, g17873)
g25940(1) = OR(g24415, g22218)
g25801(1) = AND(g8097, g24585)
g18538(1) = AND(g2759, g15277)
g24674(1) = AND(g446, g23496)
g18241(1) = AND(g1183, g16431)
g18771(1) = AND(g5685, g15615)
g18235(1) = AND(g1141, g16326)
g18683(1) = AND(g4674, g15885)
g18515(1) = AND(g2643, g15509)
g18414(1) = AND(g2102, g15373)
g18407(1) = AND(g2016, g15373)
g26085(1) = AND(g11906, g25070)
g18441(1) = AND(g2246, g18008)
g18584(1) = AND(g2950, g16349)
g18206(1) = AND(g918, g15938)
g18759(1) = AND(g5467, g17929)
g18725(1) = AND(g4912, g16077)
g25876(1) = AND(g3470, g24667)
g18114(1) = AND(g452, g17015)
g18758(1) = AND(g7004, g15595)
g24746(1) = OR(g22588, g19461)
g18435(1) = AND(g2173, g18008)
g18107(1) = AND(g429, g17015)
g18744(1) = AND(g5124, g17847)
g18345(1) = AND(g1736, g17955)
g18399(1) = AND(g2024, g15373)
g18398(1) = AND(g2020, g15373)
g18141(1) = AND(g568, g17533)
g18652(1) = AND(g4172, g16249)
g18804(1) = AND(g15163, g15656)
g18263(1) = AND(g1249, g16000)
g18332(1) = AND(g1677, g17873)
g18135(1) = AND(g136, g17249)
g18406(1) = AND(g2060, g15373)
g18361(1) = AND(g1821, g17955)
g18500(1) = AND(g2421, g15426)
g23475(1) = AND(g19070, g8971)
g18221(1) = AND(g1018, g16100)
g26815(1) = AND(g4108, g24528)
g24141(1) = AND(g17657, g21656)
g18613(1) = AND(g3338, g17200)
g18106(1) = AND(g411, g17015)
g18605(1) = AND(g3129, g16987)
g18812(1) = AND(g6509, g15483)
g18463(1) = AND(g2375, g15224)
g24406(1) = AND(g13623, g22860)
g25502(1) = AND(g6946, g22527)
g18371(1) = AND(g1870, g15171)
g18234(1) = AND(g1129, g16326)
g18795(1) = AND(g6163, g15348)
g18514(1) = AND(g2629, g15509)
g18507(1) = AND(g2595, g15509)
g25815(1) = AND(g8155, g24603)
g18163(1) = AND(g79, g17433)
g25975(1) = AND(g9434, g24999)
g18541(1) = AND(g2767, g15277)
g18473(1) = AND(g2342, g15224)
g18789(1) = AND(g6035, g15634)
g18788(1) = AND(g6031, g15634)
g18724(1) = AND(g4907, g16077)
g25884(1) = AND(g11153, g24711)
g18359(1) = AND(g1825, g17955)
g18325(1) = AND(g1624, g17873)
g18535(1) = AND(g2741, g15277)
g18434(1) = AND(g2217, g18008)
g18358(1) = AND(g1811, g17955)
g18121(1) = AND(g424, g17015)
g18344(1) = AND(g1740, g17955)
g18682(1) = AND(g4646, g15885)
g18291(1) = AND(g1437, g16449)
g18173(1) = AND(g736, g17328)
g18760(1) = AND(g5462, g17929)
g18134(1) = AND(g534, g17249)
g24959(1) = NOR(g8858, g23324)
g24724(1) = AND(g17624, g22432)
g18506(1) = AND(g2571, g15509)
g18649(1) = AND(g4049, g17271)
g18240(1) = AND(g15066, g16431)
g18648(1) = AND(g4045, g17271)
g18491(1) = AND(g2518, g15426)
g18604(1) = AND(g3125, g16987)
g18755(1) = AND(g5343, g15595)
g18770(1) = AND(g15153, g15615)
g18563(1) = AND(g2890, g16349)
g18767(1) = AND(g15150, g17929)
g18794(1) = AND(g6154, g15348)
g18395(1) = AND(g12849, g15373)
g18262(1) = AND(g1259, g16000)
g18633(1) = AND(g6905, g17226)
g18191(1) = AND(g827, g17821)
g18719(1) = AND(g4894, g16795)
g18718(1) = AND(g4854, g15915)
g18521(1) = AND(g2667, g15509)
g18440(1) = AND(g2255, g18008)
g18573(1) = AND(g2898, g16349)
g18247(1) = AND(g1178, g16431)
g23553(1) = AND(g19413, g11875)
g18389(1) = AND(g1974, g15171)
g18612(1) = AND(g3329, g17200)
g18388(1) = AND(g1968, g15171)
g18324(1) = AND(g1644, g17873)
g18701(1) = AND(g4771, g16856)
g25407(1) = NOR(g23871, g14645)
g18777(1) = AND(g5808, g18065)
g18534(1) = AND(g2735, g15277)
g18251(1) = AND(g996, g16897)
g18272(1) = AND(g1283, g16031)
g24719(1) = AND(g681, g23530)
g18462(1) = AND(g2361, g15224)
g18140(1) = AND(g559, g17533)
g26165(1) = AND(g11980, g25153)
g18766(1) = AND(g5495, g17929)
g24573(1) = AND(g17198, g23716)
g18360(1) = AND(g1830, g17955)
g18447(1) = AND(g2208, g18008)
g18162(1) = AND(g686, g17433)
g18629(1) = AND(g3680, g17226)
g18451(1) = AND(g2295, g15224)
g18472(1) = AND(g2413, g15224)
g18220(1) = AND(g1002, g16100)
g18628(1) = AND(g15095, g17226)
g24140(1) = AND(g17663, g21654)
g18246(1) = AND(g1199, g16431)
g18591(1) = AND(g2965, g16349)
g18776(1) = AND(g5813, g18065)
g18785(1) = AND(g5849, g18065)
g18147(1) = AND(g599, g17533)
g18754(1) = AND(g5339, g15595)
g18355(1) = AND(g1748, g17955)
g18825(1) = AND(g6736, g15680)
g18370(1) = AND(g1874, g15171)
g18151(1) = AND(g617, g17533)
g18172(1) = AND(g15058, g17328)
g18367(1) = AND(g1783, g17955)
g18394(1) = AND(g1862, g15171)
g26021(1) = AND(g9568, g25035)
g18420(1) = AND(g1996, g15373)
g18319(1) = AND(g1600, g17873)
g18318(1) = AND(g1604, g17873)
g18446(1) = AND(g2279, g18008)
g18227(1) = AND(g1052, g16129)
g18540(1) = AND(g2775, g15277)
g25063(1) = AND(g13078, g22325)
g18203(1) = AND(g911, g15938)
g18281(1) = AND(g1373, g16136)
g18301(1) = AND(g1532, g16489)
g18377(1) = AND(g1894, g15171)
g18120(1) = AND(g457, g17015)
g18739(1) = AND(g5008, g16826)
g18146(1) = AND(g595, g17533)
g18738(1) = AND(g15142, g16826)
g18645(1) = AND(g15100, g17271)
g23997(1) = OR(g20602, g17191)
g25321(1) = NOR(g23835, g14645)
g18699(1) = AND(g4760, g16816)
g18290(1) = AND(g1467, g16449)
g18698(1) = AND(g15131, g16777)
g18427(1) = AND(g2181, g18008)
g18366(1) = AND(g1854, g17955)
g18632(1) = AND(g3698, g17226)
g25446(1) = NOR(g23686, g14645)
g18403(1) = AND(g2028, g15373)
g18547(1) = AND(g121, g15277)
g25565(1) = AND(g13013, g22660)
g18226(1) = AND(g15064, g16129)
g18715(1) = AND(g4871, g15915)
g18481(1) = AND(g2461, g15426)
g18551(1) = AND(g2811, g15277)
g18572(1) = AND(g2864, g16349)
g18127(1) = AND(g499, g16971)
g18490(1) = AND(g2504, g15426)
g18784(1) = AND(g15155, g18065)
g18376(1) = AND(g1913, g15171)
g18385(1) = AND(g1959, g15171)
g18297(1) = AND(g1478, g16449)
g18103(1) = AND(g401, g17015)
g18354(1) = AND(g1792, g17955)
g18824(1) = AND(g6732, g15680)
g18181(1) = AND(g772, g17328)
g18671(1) = AND(g4628, g15758)
g23998(1) = AND(g19631, g10971)
g24551(1) = AND(g17148, g23331)
g18426(1) = AND(g2177, g18008)
g18190(1) = AND(g822, g17821)
g23513(1) = AND(g19430, g13007)
g18520(1) = AND(g2661, g15509)
g18546(1) = AND(g2795, g15277)
g18211(1) = AND(g15062, g15979)
g18497(1) = AND(g2541, g15426)
g18700(1) = AND(g15132, g16816)
g18126(1) = AND(g15054, g16971)
g18659(1) = AND(g4366, g17183)
g18625(1) = AND(g15092, g17062)
g18250(1) = AND(g6821, g16897)
g18658(1) = AND(g15121, g17183)
g25522(1) = AND(g6888, g22544)
g18339(1) = AND(g1714, g17873)
g18296(1) = AND(g1495, g16449)
g18644(1) = AND(g15098, g17125)
g18338(1) = AND(g1710, g17873)
g22447(1) = OR(g21464, g12761)
g18197(1) = AND(g854, g17821)
g18411(1) = AND(g2093, g15373)
g24700(1) = AND(g645, g23512)
g18503(1) = AND(g2563, g15509)
g18581(1) = AND(g2912, g16349)
g18714(1) = AND(g4864, g15915)
g24896(1) = OR(g22863, g19684)
g18450(1) = AND(g2299, g15224)
g18315(1) = AND(g1548, g16931)
g18707(1) = AND(g15134, g16782)
g18819(1) = AND(g6541, g15483)
g18202(1) = AND(g907, g15938)
g18257(1) = AND(g1205, g16897)
g26780(1) = AND(g4098, g24437)
g18818(1) = AND(g15165, g15483)
g18496(1) = AND(g2537, g15426)
g18111(1) = AND(g174, g17015)
g25872(1) = AND(g3119, g24655)
g18590(1) = AND(g2917, g16349)
g18741(1) = AND(g15143, g17384)
g18384(1) = AND(g1945, g15171)
g18150(1) = AND(g604, g17533)
g18801(1) = AND(g15160, g15348)
g18735(1) = AND(g4983, g16826)
g18196(1) = AND(g703, g17821)
g18526(1) = AND(g2555, g15509)
g25943(1) = OR(g24423, g22299)
g26020(1) = AND(g9559, g25034)
g25942(1) = OR(g24422, g22298)
g18402(1) = AND(g2047, g15373)
g18457(1) = AND(g2319, g15224)
g18706(1) = AND(g4785, g16782)
g25834(1) = OR(g25366, g23854)
g18256(1) = AND(g1242, g16897)
g18689(1) = AND(g15129, g16752)
g18280(1) = AND(g1367, g16136)
g18688(1) = AND(g4704, g16752)
g18624(1) = AND(g3490, g17062)
g18300(1) = AND(g1306, g16489)
g23533(1) = AND(g19436, g13015)
g18157(1) = AND(g15057, g17433)
g18231(1) = AND(g1105, g16326)
g25022(1) = NOR(g714, g23324)
g24001(1) = AND(g19651, g10951)
g18511(1) = AND(g2599, g15509)
g18763(1) = AND(g5481, g17929)
g21512(1) = AND(g16225, g10881)
g18456(1) = AND(g2338, g15224)
g25501(1) = NOR(g23918, g14645)
g18480(1) = AND(g2437, g15426)
g20271(1) = NAND(g16925, g14054, g16657, g16628)
g20150(1) = NAND(g17705, g17669, g17635, g14590)
g21555(1) = NAND(g17846, g14946, g17686, g17650)
g21364(1) = NAND(g15787, g15781, g15753, g13131)
g21603(1) = NAND(g17872, g14987, g17723, g17689)
g21386(1) = NAND(g15798, g15788, g15782, g13139)
g20371(1) = NAND(g16956, g14088, g16694, g16660)
g20161(1) = NAND(g17732, g17706, g17670, g14625)
g21509(1) = NAND(g17820, g14898, g17647, g17608)
g21356(1) = NAND(g15780, g15752, g15743, g13118)
g21429(1) = NAND(g17788, g14803, g17578, g17520)
g21338(1) = NAND(g15741, g15734, g15728, g13097)
g20236(1) = NAND(g16875, g14014, g16625, g16604)
g20133(1) = NAND(g17668, g17634, g17597, g14569)
g21459(1) = NAND(g17814, g14854, g17605, g17581)
g21350(1) = NAND(g15751, g15742, g15735, g13108)
I20165(2) = NAND(g16246, g990)
I20221(2) = NAND(g16272, g11170)
g22642(1) = NAND(g7870, g19560)
I23118(2) = NAND(g20076, g417)
g23379(1) = NAND(g20216, g11248)
I20203(2) = NAND(g16246, g11147)
g22833(1) = NAND(g1193, g19560, g10666)
g26752(1) = NAND(g9397, g25189)
g26255(1) = NAND(g8075, g24779)
g26782(1) = NAND(g9467, g25203)
g22687(1) = NAND(g19560, g7870)
g22711(1) = NAND(g19581, g7888)
I16780(1) = NAND(g12332, I16778)
I16779(1) = NAND(g11292, I16778)
g26235(1) = NAND(g8016, g24766)
I20187(2) = NAND(g16272, g1333)
g26208(1) = NAND(g7975, g24751)
g26714(1) = NAND(g9316, g25175)
g26685(1) = NAND(g9264, g25160)
g22850(1) = NAND(g1536, g19581, g10699)
g22650(1) = NAND(g7888, g19581)
g26666(1) = NAND(g9229, g25144)
g23357(1) = NAND(g20201, g11231)
g23190(1) = NOT(I22286)
g24151(1) = OR(g18088, g21661)
I21294(1) = NOT(g18274)
g20785(52) = NOT(I20846)
g24066(1) = NOT(g21127)
I22692(1) = NOT(g21308)
g19801(50) = NOT(I20216)
g21611(40) = NOT(I21210)
I21285(1) = NOT(g18215)
I22400(1) = NOT(g19620)
g18833(40) = NOT(I19661)
g27015(1) = NOT(g26869)
g19277(52) = NOT(I19813)
g18997(52) = NOT(I19756)
g26672(1) = NOT(g25275)
I20816(1) = NOT(g17088)
g21514(40) = NOT(I21189)
I21002(1) = NOT(g16709)
g19074(52) = NOT(I19772)
I22539(1) = NOT(g19606)
g19210(52) = NOT(I19796)
I21776(1) = NOT(g21308)
g19147(52) = NOT(I19786)
g24076(1) = NOT(g19984)
g24085(1) = NOT(g20857)
g20596(1) = NOT(I20690)
g23764(2) = NOT(g21308)
g24054(1) = NOT(g19919)
g27295(2) = NAND(g24776, g26208)
I20753(1) = NOT(g16677)
I23312(1) = NOT(g21681)
g21070(52) = NOT(I20937)
g20924(52) = NOT(I20895)
I22343(1) = NOT(g19371)
g24131(1) = NOT(g21209)
I20233(1) = NOT(g17487)
I21477(1) = NOT(g18695)
I20647(1) = NOT(g17010)
I22114(1) = NOT(g19935)
g21468(40) = NOT(I21181)
g27242(1) = NOT(g26183)
g24039(1) = NOT(g21256)
g24038(1) = NOT(g21193)
I22583(1) = NOT(g20998)
I21036(1) = NOT(g17221)
g20453(40) = NOT(I20584)
g21562(40) = NOT(I21199)
I22561(1) = NOT(g20841)
g20283(36) = NOT(I20529)
g26681(1) = NOT(g25396)
g25888(3) = NAND(g914, g24439)
I22425(1) = NOT(g19379)
g23828(6) = AND(g9104, g19128)
g26765(1) = NOT(g25309)
g20391(40) = NOT(I20562)
g27237(1) = NOT(g26162)
g24084(1) = NOT(g20720)
g24110(1) = NOT(g21209)
I21941(1) = NOT(g18918)
g22908(10) = NAND(g9104, g20175)
I20750(1) = NOT(g16677)
I22622(1) = NOT(g21209)
g23816(2) = NOT(g21308)
g24964(1) = NOT(I24128)
g22138(1) = NOT(g21370)
I20982(1) = NOT(g16300)
g18940(2) = NOT(I19719)
g24117(1) = NOT(g21209)
g22942(14) = AND(g9104, g20219)
g24123(1) = NOT(g21143)
g23865(2) = NOT(g21308)
I22028(1) = NOT(g20204)
g26736(1) = NOT(g25349)
g20330(40) = NOT(I20542)
I20999(1) = NOT(g16709)
g23267(2) = NOT(g20097)
I22240(1) = NOT(g20086)
I22604(1) = NOT(g21143)
g23742(2) = AND(g19128, g9104)
g24116(1) = NOT(g21143)
I22316(1) = NOT(g19361)
g26709(1) = NOT(g25435)
g27565(1) = NOT(g26645)
g24041(1) = NOT(g19968)
I21787(1) = NOT(g19422)
g24035(1) = NOT(g20841)
g21273(1) = NOT(I21006)
I22380(1) = NOT(g21156)
I22619(1) = NOT(g21193)
I22000(1) = NOT(g20277)
g21037(10) = NOT(I20913)
g24130(1) = NOT(g20998)
g26792(1) = NOT(g25439)
g23802(6) = AND(g9104, g19050)
g27670(2) = NAND(g25172, g26666)
g26598(3) = NOR(g8990, g13756, g24732)
g22885(10) = NAND(g9104, g20154)
g24575(1) = NOR(g23498, g23514)
g24063(1) = NOT(g20014)
g26656(1) = NOT(g25495)
g24137(1) = NOT(g20998)
g22670(8) = AND(g20114, g9104)
g26680(1) = NOT(g25300)
g27020(3) = AND(g4601, g25852)
I20957(1) = NOT(g16228)
g26631(1) = NOT(g25467)
I21838(1) = NOT(g19263)
g24021(1) = NOT(g20841)
g24073(1) = NOT(g21127)
I21744(1) = NOT(g19338)
I21849(1) = NOT(g19620)
g24122(1) = NOT(g20857)
g24034(1) = NOT(g19968)
I23303(1) = NOT(g21669)
g24136(1) = NOT(g20857)
g23239(2) = NOT(g21308)
g27629(3) = NOR(g8891, g26382, g12259)
I20954(1) = NOT(g16228)
I22264(1) = NOT(g20100)
g27592(1) = NOT(g26715)
g24109(1) = NOT(g21143)
g24108(1) = NOT(g20998)
I21911(1) = NOT(g21278)
I21033(1) = NOT(g17221)
g26679(1) = NOT(g25385)
I22366(1) = NOT(g19757)
g24091(1) = NOT(g20720)
I22547(1) = NOT(g20720)
g22682(1) = NOT(g19379)
I21757(1) = NOT(g21308)
g27583(1) = NOT(g26686)
g22689(8) = AND(g18918, g9104)
g18926(2) = NOT(I19707)
g24040(1) = NOT(g19919)
I22128(1) = NOT(g19968)
I21291(1) = NOT(g18273)
g24062(1) = NOT(g19968)
I22211(1) = NOT(g21463)
g24047(1) = NOT(g19919)
g24051(1) = NOT(g21127)
g24072(1) = NOT(g20982)
I23300(1) = NOT(g21665)
g19458(2) = NOT(I19927)
g26693(1) = NOT(g25300)
I22111(1) = NOT(g19919)
g24020(1) = NOT(g20014)
g27693(2) = NAND(g25216, g26752)
I19671(1) = NOT(g15932)
g24046(1) = NOT(g21256)
I22525(1) = NOT(g19345)
I23324(1) = NOT(g21697)
g24113(1) = NOT(g19984)
I21802(1) = NOT(g21308)
g24105(1) = NOT(g19935)
g27687(2) = NAND(g25200, g26714)
I21766(1) = NOT(g19620)
I21734(1) = NOT(g19268)
g24027(1) = NOT(g20014)
I20650(1) = NOT(g17010)
I21831(1) = NOT(g19127)
g24081(1) = NOT(g21209)
I22464(1) = NOT(g21222)
g26284(1) = NOT(g24875)
g24090(1) = NOT(g19935)
I22143(1) = NOT(g20189)
g26653(1) = NOT(g25337)
I22009(1) = NOT(g21269)
I23318(1) = NOT(g21689)
g24026(1) = NOT(g19919)
g27245(1) = NOT(g26209)
g24149(1) = NOT(g19338)
g21366(2) = NOT(I21100)
g24097(1) = NOT(g19935)
g24104(1) = NOT(g19890)
I22131(1) = NOT(g19984)
g23789(2) = NOT(g21308)
I22458(1) = NOT(g18954)
I22502(1) = NOT(g19376)
I22153(1) = NOT(g20014)
g20695(1) = NOT(I20781)
I19674(1) = NOT(g15932)
g24133(1) = NOT(g19935)
g26732(1) = NOT(g25389)
I22601(1) = NOT(g21127)
I21918(1) = NOT(g21290)
I20321(1) = NOT(g16920)
g24112(1) = NOT(g19935)
g24050(1) = NOT(g20841)
I21784(1) = NOT(g19638)
I21297(1) = NOT(g18597)
g24096(1) = NOT(g19890)
I21969(1) = NOT(g21370)
g26683(1) = NOT(g25514)
I21480(1) = NOT(g18696)
I22580(1) = NOT(g20982)
g23599(2) = AND(g19050, g9104)
I20985(1) = NOT(g16300)
I21860(1) = NOT(g19638)
g24129(1) = NOT(g20857)
g24057(1) = NOT(g20841)
g24128(1) = NOT(g20720)
g23191(1) = NOT(I22289)
g22876(4) = AND(g20136, g9104)
g22714(1) = NOT(g20436)
I24558(1) = NOT(g23777)
g26758(1) = NOT(g25389)
g26744(1) = NOT(g25400)
g26804(1) = NOT(g25400)
I22665(1) = NOT(g21308)
g22150(1) = NOT(g21280)
I22589(1) = NOT(g21340)
I23315(1) = NOT(g21685)
g24056(1) = NOT(g20014)
g24080(1) = NOT(g21143)
I22461(1) = NOT(g21225)
g24031(1) = NOT(g21193)
I22124(1) = NOT(g21300)
I21815(1) = NOT(g21308)
g26812(1) = NOT(g25439)
I21019(1) = NOT(g17325)
g25895(3) = NAND(g1259, g24453)
I20819(1) = NOT(g17088)
g24132(1) = NOT(g19890)
I22275(1) = NOT(g20127)
I22046(1) = NOT(g19330)
g24087(1) = NOT(g21143)
g23844(2) = NOT(g21308)
I22499(1) = NOT(g21160)
g24043(1) = NOT(g20982)
I21300(1) = NOT(g18598)
g24069(1) = NOT(g19968)
g26788(1) = NOT(g25349)
g26724(1) = NOT(g25341)
g24068(1) = NOT(g19919)
I20864(1) = NOT(g16960)
g26682(1) = NOT(g25309)
g24079(1) = NOT(g20998)
g18562(1) = NOT(I19384)
g22667(1) = NOT(g21156)
g24078(1) = NOT(g20857)
g24086(1) = NOT(g20998)
I22542(1) = NOT(g19773)
I21792(1) = NOT(g21308)
I20867(1) = NOT(g16216)
I23321(1) = NOT(g21693)
g24125(1) = NOT(g19890)
I22512(1) = NOT(g19389)
I21930(1) = NOT(g21297)
I22422(1) = NOT(g19330)
I22488(1) = NOT(g18984)
g27306(2) = NAND(g24787, g26235)
g24023(1) = NOT(g21127)
g26820(1) = NOT(I25534)
I23306(1) = NOT(g21673)
g23211(2) = NOT(g21308)
g26701(1) = NOT(g25341)
g26777(1) = NOT(g25439)
I21486(1) = NOT(g18727)
I22327(1) = NOT(g19367)
g21335(1) = NOT(I21067)
g24042(1) = NOT(g20014)
g24124(1) = NOT(g21209)
g23639(2) = AND(g19050, g9104)
g24030(1) = NOT(g21127)
g24093(1) = NOT(g20998)
g26776(1) = NOT(g25498)
I22571(1) = NOT(g20097)
g24065(1) = NOT(g20982)
g26754(1) = NOT(g25300)
g25766(1) = NOT(g24439)
I22302(1) = NOT(g19353)
I22485(1) = NOT(g21308)
g27317(2) = NAND(g24793, g26255)
I22564(1) = NOT(g20857)
g24075(1) = NOT(g19935)
g23076(2) = AND(g19128, g9104)
g24037(1) = NOT(g21127)
I23309(1) = NOT(g21677)
g26632(1) = NOT(g25473)
g24119(1) = NOT(g19935)
g26352(3) = NAND(g744, g24875, g11679)
g24118(1) = NOT(g19890)
g24022(1) = NOT(g20982)
g23675(2) = AND(g19050, g9104)
I22640(1) = NOT(g21256)
g24053(1) = NOT(g21256)
g24036(1) = NOT(g20982)
g24101(1) = NOT(g20998)
g27415(1) = NOT(g26382)
g26784(1) = NOT(g25341)
g24064(1) = NOT(g20841)
I20744(1) = NOT(g17141)
g27554(1) = NOT(g26625)
g22137(1) = NOT(g21370)
g24074(1) = NOT(g21193)
g26700(1) = NOT(g25429)
g24092(1) = NOT(g20857)
g22136(1) = NOT(g20277)
g24083(1) = NOT(g19984)
I22470(1) = NOT(g21326)
I22331(1) = NOT(g19417)
I20747(1) = NOT(g17141)
g27991(1) = NOT(g25852)
g23708(2) = AND(g19050, g9104)
g23223(2) = NOT(g21308)
g23958(2) = AND(g9104, g19200)
g24138(1) = NOT(g21143)
g23121(2) = AND(g19128, g9104)
I22149(1) = NOT(g21036)
g24115(1) = NOT(g20998)
g27965(1) = AND(g25834, g13117)
g24052(1) = NOT(g21193)
I21483(1) = NOT(g18726)
I22096(1) = NOT(g19890)
g19699(9) = NOT(I20116)
g24100(1) = NOT(g20857)
I20861(1) = NOT(g16960)
g22756(1) = NOT(g20436)
g26655(1) = NOT(g25492)
g24114(1) = NOT(g20720)
g24082(1) = NOT(g19890)
g24107(1) = NOT(g20857)
I22467(1) = NOT(g19662)
g25773(1) = NOT(g24453)
g25930(1) = NOT(I25028)
I22444(1) = NOT(g19626)
g24135(1) = NOT(g20720)
g21175(1) = NOT(I20951)
I20318(1) = NOT(g16920)
g24049(1) = NOT(g20014)
g24048(1) = NOT(g19968)
g21387(1) = NOT(I21115)
g24106(1) = NOT(g19984)
I21769(1) = NOT(g19402)
g24033(1) = NOT(g19919)
I21959(1) = NOT(g20242)
g26654(1) = NOT(g25275)
g25222(1) = NOT(I24400)
I22419(1) = NOT(g19638)
g27573(1) = NOT(g26667)
g24121(1) = NOT(g20720)
g22646(1) = NOT(g19389)
g24134(1) = NOT(g19984)
g24029(1) = NOT(g20982)
I25750(1) = NOT(g26823)
g24506(1) = NOT(I23711)
g24028(1) = NOT(g20841)
I22353(1) = NOT(g19375)
g23148(2) = AND(g19128, g9104)
g26615(1) = NOT(g25432)
g26720(1) = NOT(g25275)
g23314(2) = AND(g9104, g19200)
g27679(2) = NAND(g25186, g26685)
g24045(1) = NOT(g21193)
I20870(1) = NOT(g16216)
g24099(1) = NOT(g20720)
g24098(1) = NOT(g19984)
g24032(1) = NOT(g21256)
g24061(1) = NOT(g19919)
g24071(1) = NOT(g20841)
g26614(1) = NOT(g25426)
g24147(1) = NOT(g19402)
g26607(1) = NOT(g25382)
g24059(1) = NOT(g21193)
g24025(1) = NOT(g21256)
g24058(1) = NOT(g20982)
g24044(1) = NOT(g21127)
g24120(1) = NOT(g19984)
g24146(1) = NOT(g19422)
g22994(1) = NOT(g20436)
g24127(1) = NOT(g19984)
g24103(1) = NOT(g21209)
g24095(1) = NOT(g21209)
g26702(1) = NOT(g25309)
I21288(1) = NOT(g18216)
g26634(1) = NOT(g25317)
g19720(9) = NOT(I20130)
g24089(1) = NOT(g19890)
g26745(3) = NAND(g6856, g25317)
g24088(1) = NOT(g21209)
g24024(1) = NOT(g21193)
g24126(1) = NOT(g19935)
I22729(1) = NOT(g21308)
g24060(1) = NOT(g21256)
g26731(1) = NOT(g25470)
g23293(2) = AND(g9104, g19200)
g24055(1) = NOT(g19968)
g24111(1) = NOT(g19890)
g24070(1) = NOT(g20014)
g24067(1) = NOT(g21256)
g24094(1) = NOT(g21143)
g26743(1) = NOT(g25476)
g24150(1) = NOT(g19268)
g24019(1) = NOT(g19968)
g26769(1) = NOT(g25400)
g26803(1) = NOT(g25389)
g26330(3) = NOR(g8631, g24825)
g27038(1) = NOT(g25932)
g24077(1) = NOT(g20720)
g26710(1) = NOT(g25349)
g27705(2) = NAND(g25237, g26782)
g24619(1) = NOR(g23554, g23581)
g24102(1) = NOT(g21143)
g22623(1) = AND(g19337, g19470)
g24907(1) = OR(g21558, g24015)
g23056(1) = AND(g16052, g19860)
g26090(1) = AND(g1624, g25081)
g26233(1) = AND(g2279, g25309)
g26182(1) = AND(g9978, g25317)
g24660(1) = AND(g22648, g19737)
g22589(1) = AND(g19267, g19451)
g27574(1) = OR(g26145, g24730)
g26377(1) = OR(g24700, g23007)
g24773(1) = AND(g22832, g19872)
g26387(1) = AND(g24813, g20231)
g23471(1) = AND(g20148, g20523)
g26104(1) = AND(g2250, g25101)
g22900(1) = AND(g17137, g19697)
g26309(1) = NOR(g8575, g24825)
g27533(1) = OR(g26078, g24659)
g23774(1) = AND(g14867, g21252)
g22929(5) = NOR(g19773, g12970)
g24502(1) = AND(g23428, g13223)
g24618(1) = AND(g22625, g19672)
g26229(1) = AND(g1724, g25275)
g26310(1) = AND(g2102, g25389)
g25906(1) = OR(g25559, g24014)
g25971(1) = AND(g1917, g24992)
g23901(1) = AND(g19606, g7963)
g22518(1) = AND(g12982, g19398)
g22637(1) = AND(g19363, g19489)
g27275(1) = AND(g25945, g19745)
g25959(1) = AND(g1648, g24963)
g26346(1) = NOR(g8522, g24825)
g25925(1) = AND(g24990, g23234)
g26129(1) = AND(g2384, g25121)
g26386(1) = OR(g24719, g23023)
g27555(1) = OR(g26095, g24686)
g26128(1) = AND(g2319, g25120)
g27544(1) = OR(g26087, g24671)
g22622(1) = AND(g19336, g19469)
g26232(1) = AND(g2193, g25396)
g27429(1) = OR(g25969, g24589)
g27456(1) = OR(g25978, g24607)
g25057(1) = AND(g23275, g20511)
g27133(1) = OR(g25788, g24392)
g27821(1) = AND(g7680, g25892)
g26611(1) = AND(g24935, g20580)
g27264(1) = AND(g25941, g19714)
g26271(1) = AND(g1992, g25341)
g23188(1) = AND(g13994, g20025)
g27226(1) = OR(g25872, g24436)
g26161(1) = AND(g2518, g25139)
g25924(1) = AND(g24976, g16846)
g23218(1) = AND(g20200, g16530)
g22329(1) = AND(g11940, g20329)
g23837(1) = AND(g21160, g10804)
g24983(1) = AND(g23217, g20238)
g27239(1) = OR(g25881, g24465)
g26602(1) = AND(g7487, g24453)
g23201(1) = AND(g14027, g20040)
g27426(1) = OR(g25967, g24588)
g24523(1) = AND(g22318, g19468)
g22515(1) = AND(g12981, g19395)
g25069(1) = AND(g23296, g20535)
g25955(1) = AND(g24720, g19580)
g24600(1) = AND(g22591, g19652)
g25970(1) = AND(g1792, g24991)
g26159(1) = AND(g2370, g25137)
g26125(1) = AND(g1894, g25117)
g26158(1) = AND(g2255, g25432)
g26783(1) = AND(g25037, g21048)
g22849(1) = AND(g1227, g19653)
g23254(1) = AND(g20056, g20110)
g22848(1) = AND(g19449, g19649)
g25078(1) = AND(g23298, g20538)
g26289(1) = AND(g2551, g25400)
g24853(1) = OR(g21452, g24001)
g26288(1) = AND(g2259, g25309)
g23166(1) = AND(g13959, g19979)
g23008(1) = AND(g1570, g19783)
g24797(1) = AND(g22872, g19960)
g24408(1) = AND(g23989, g18946)
g26544(1) = AND(g7446, g24357)
g26713(1) = AND(g25447, g20714)
g27820(1) = AND(g7670, g25932)
g23439(1) = AND(g13771, g20452)
g26270(1) = AND(g1700, g25275)
g26124(1) = AND(g1811, g25116)
g23349(1) = AND(g13662, g20182)
g23083(1) = AND(g16076, g19878)
g25545(1) = OR(g23551, g20658)
g24553(1) = AND(g22983, g19539)
g26160(1) = AND(g2453, g25138)
g23415(1) = AND(g20077, g20320)
g25042(1) = AND(g23262, g20496)
g26972(1) = OR(g26780, g25229)
g24583(1) = NAND(g22753, g22711)
g26277(1) = AND(g2547, g25400)
g25030(1) = AND(g23251, g20432)
g23484(1) = AND(g20160, g20541)
g24673(1) = AND(g22659, g19748)
g26155(1) = AND(g1945, g25134)
g24841(1) = OR(g21420, g23998)
g23921(1) = AND(g19379, g4146)
g24634(1) = AND(g22634, g19685)
g27249(1) = AND(g25929, g19678)
g23799(1) = AND(g14911, g21279)
g27403(1) = OR(g25962, g24581)
g26422(1) = OR(g24774, g23104)
g22899(1) = AND(g19486, g19695)
g22990(1) = AND(g19555, g19760)
g24926(2) = NAND(g20172, g20163, g23357, g13995)
g22633(1) = AND(g19359, g19479)
g24494(1) = NOR(g23513, g23532)
g26276(1) = AND(g2461, g25476)
g26285(1) = AND(g1834, g25300)
g26254(1) = AND(g2413, g25349)
g26808(1) = AND(g25521, g21185)
g26101(1) = AND(g1760, g25098)
g26177(1) = AND(g2079, g25154)
g26512(1) = OR(g24786, g23130)
g23991(1) = AND(g19209, g21428)
g25867(1) = OR(g25449, g23884)
g25900(1) = AND(g24390, g19368)
g23407(1) = AND(g9295, g20273)
g25466(1) = AND(g23574, g21346)
g24508(1) = NOR(g23577, g23618)
g24743(1) = AND(g22708, g19789)
g24803(1) = AND(g22901, g20005)
g23725(1) = AND(g14772, g21138)
g26176(1) = AND(g1964, g25467)
g26092(1) = AND(g9766, g25083)
g26154(1) = AND(g1830, g25426)
g27147(1) = OR(g25802, g24399)
g27524(1) = OR(g26050, g24649)
g24710(1) = AND(g22679, g19771)
g27378(1) = AND(g26089, g20052)
g22487(1) = OR(g21512, g12794)
g24945(1) = AND(g23183, g20197)
g26267(1) = NOR(g8033, g24732)
g25883(1) = AND(g13728, g24699)
g26247(1) = NOR(g7995, g24732)
g24961(1) = AND(g23193, g20209)
g24717(1) = AND(g22684, g19777)
g22632(1) = AND(g19356, g19476)
g26268(1) = NOR(g283, g24825)
g24646(1) = AND(g22640, g19711)
g26799(1) = AND(g25247, g21068)
g23724(1) = AND(g14767, g21123)
g25963(1) = AND(g1657, g24978)
g27233(1) = OR(g25876, g24451)
g23682(1) = AND(g16970, g20874)
g24936(2) = NAND(g20186, g20173, g23379, g14029)
g26207(1) = AND(g2638, g25170)
g27556(1) = OR(g26097, g24687)
g27145(1) = AND(g14121, g26382)
g25973(1) = AND(g2342, g24994)
g26100(1) = AND(g1677, g25097)
g23755(1) = AND(g14821, g21204)
g24504(1) = AND(g22226, g19410)
g26206(1) = AND(g2523, g25495)
g22590(1) = AND(g19274, g19452)
g25991(1) = AND(g2060, g25023)
g23389(1) = AND(g9072, g19757)
g25836(1) = OR(g25368, g23856)
g24499(1) = AND(g22217, g19394)
g26609(1) = NOR(g146, g24732)
g25539(1) = OR(g23531, g20628)
g26273(1) = AND(g2122, g25389)
g23451(1) = AND(g13805, g20510)
g24650(1) = AND(g22641, g19718)
g23220(1) = AND(g19417, g20067)
g22624(1) = AND(g19344, g19471)
g26234(1) = AND(g2657, g25514)
g22157(1) = AND(g14608, g18892)
g23754(1) = AND(g14816, g21189)
g27232(1) = OR(g25874, g24450)
g26514(1) = AND(g7400, g25564)
g27179(1) = OR(g25816, g24409)
g25951(1) = AND(g24500, g19565)
g25972(1) = AND(g2217, g24993)
g24657(1) = AND(g22644, g19730)
g23025(1) = AND(g16021, g19798)
g24919(1) = OR(g21606, g22143)
g23540(1) = AND(g16866, g20622)
g24967(1) = AND(g23197, g20213)
g26291(1) = AND(g2681, g25439)
g27584(1) = OR(g26165, g24758)
g27575(1) = OR(g26147, g24731)
g27255(1) = AND(g25936, g19689)
g25946(1) = AND(g24496, g19537)
g24532(1) = AND(g22331, g19478)
g24977(1) = AND(g23209, g20232)
g23572(1) = AND(g20230, g20656)
g27160(1) = AND(g14163, g26340)
g26845(1) = AND(g24391, g21426)
g26359(1) = OR(g24651, g22939)
g25927(1) = AND(g25004, g20375)
g27205(1) = OR(g25833, g24421)
g25491(1) = AND(g23615, g21355)
g25981(1) = AND(g2051, g25007)
g26324(1) = AND(g2661, g25439)
g26251(1) = AND(g1988, g25341)
g24643(1) = AND(g22636, g19696)
g26272(1) = AND(g2036, g25470)
g23497(1) = AND(g20169, g20569)
g24669(1) = AND(g22653, g19742)
g26338(1) = NOR(g8458, g24825)
g25877(1) = OR(g25502, g23919)
g23658(1) = AND(g14687, g20852)
g24559(1) = AND(g22993, g19567)
g24016(1) = AND(g14528, g21610)
g22516(1) = OR(g21559, g12817)
g26349(1) = OR(g24630, g13409)
g25926(1) = AND(g25005, g24839)
g27254(1) = AND(g25935, g19688)
g27506(1) = OR(g26021, g24639)
g26299(1) = OR(g24551, g22665)
g27567(1) = OR(g26121, g24714)
g26844(1) = AND(g25261, g21418)
g22992(1) = AND(g1227, g19765)
g24915(1) = AND(g23087, g20158)
g22835(1) = AND(g15803, g19633)
g26298(1) = NOR(g8297, g24825)
g26203(1) = AND(g1632, g25337)
g27487(1) = OR(g25990, g24629)
g26290(1) = AND(g2595, g25498)
g23280(1) = AND(g19417, g20146)
g27453(1) = OR(g25976, g24606)
g25058(1) = AND(g23276, g20513)
g25819(1) = OR(g25323, g23836)
g22165(1) = AND(g15594, g18903)
g25902(1) = AND(g24398, g19373)
g25957(1) = AND(g17190, g24960)
g26572(1) = AND(g7443, g24439)
g26127(1) = AND(g2236, g25119)
g26103(1) = AND(g2185, g25100)
g26181(1) = AND(g2652, g25157)
g27484(1) = OR(g25988, g24628)
g25551(1) = AND(g23822, g21511)
g22834(1) = AND(g102, g19630)
g26024(1) = AND(g2619, g25039)
g23131(1) = AND(g13919, g19930)
g26628(1) = NOR(g8990, g24732)
g25980(1) = AND(g1926, g25006)
g26296(1) = NOR(g8287, g24732)
g25095(1) = AND(g23319, g20556)
g24941(1) = AND(g23171, g20190)
g26126(1) = AND(g1959, g25118)
g25181(1) = AND(g23405, g20696)
g26250(1) = AND(g1902, g25429)
g26392(1) = OR(g24745, g23050)
g24574(1) = NAND(g22709, g22687)
g23187(1) = AND(g13989, g20010)
g25089(1) = AND(g23317, g20553)
g25910(1) = OR(g25565, g22142)
g22864(1) = NAND(g7780, g21156)
g24840(1) = OR(g21419, g23996)
g22982(1) = AND(g19535, g19747)
g24664(1) = AND(g22652, g19741)
g23373(1) = AND(g13699, g20195)
g24554(1) = AND(g22490, g19541)
g25979(1) = AND(g24517, g19650)
g27243(1) = OR(g25884, g24475)
g22862(1) = AND(g1570, g19673)
g25094(1) = AND(g23318, g20554)
g27263(1) = AND(g25940, g19713)
g26300(1) = AND(g1968, g25341)
g26102(1) = AND(g1825, g25099)
g26157(1) = AND(g2093, g25136)
g25526(1) = AND(g23720, g21400)
g26231(1) = AND(g1854, g25300)
g24761(1) = AND(g22751, g19852)
g22851(1) = AND(g496, g19654)
g25077(1) = AND(g23297, g20536)
g23265(1) = AND(g20069, g20132)
g23416(1) = AND(g20082, g20321)
g25923(1) = AND(g24443, g19443)
g26341(1) = AND(g24746, g20105)
g26156(1) = AND(g2028, g25135)
g27566(1) = OR(g26119, g24713)
g26180(1) = AND(g2587, g25156)
g25916(1) = AND(g24432, g19434)
g23165(1) = AND(g13954, g19964)
g26286(1) = AND(g2126, g25389)
g23006(1) = AND(g19575, g19776)
g25993(1) = AND(g2610, g25025)
g25965(1) = AND(g2208, g24980)
g24962(1) = AND(g23194, g20210)
g23372(1) = AND(g16448, g20194)
g24004(1) = AND(g37, g21225)
g23873(1) = AND(g21222, g10815)
g22710(1) = AND(g19358, g19600)
g26297(1) = NOR(g8519, g24825)
g26179(1) = AND(g2504, g25155)
g26178(1) = AND(g2389, g25473)
g24507(1) = AND(g22304, g19429)
g24012(1) = AND(g14496, g21561)
g25868(1) = OR(g25450, g23885)
g25922(1) = AND(g24959, g20065)
g25885(1) = OR(g25522, g23957)
g23474(1) = AND(g13830, g20533)
g24682(1) = AND(g22662, g19754)
g22149(1) = AND(g14581, g18880)
g26123(1) = AND(g1696, g25382)
g26230(1) = AND(g1768, g25385)
g25964(1) = AND(g1783, g24979)
g23606(1) = AND(g16927, g20679)
g27150(1) = OR(g25804, g24400)
g26098(1) = NOR(g9073, g24732)
g25909(1) = AND(g8745, g24875)
g25543(1) = AND(g23795, g21461)
g22310(1) = AND(g19662, g20235)
g26275(1) = AND(g2417, g25349)
g25992(1) = AND(g2485, g25024)
g26684(1) = AND(g25407, g20673)
g23564(1) = AND(g16882, g20648)
g23397(1) = AND(g11154, g20239)
g25041(1) = AND(g23261, g20494)
g25878(1) = OR(g25503, g23920)
g23872(1) = AND(g19389, g4157)
g26396(1) = OR(g24762, g23062)
g25983(1) = AND(g2476, g25009)
g26253(1) = AND(g2327, g25435)
g25130(1) = AND(g23358, g20600)
g24821(1) = OR(g21404, g23990)
g27543(1) = OR(g26085, g24670)
g23396(1) = AND(g20051, g20229)
g22831(1) = AND(g19441, g19629)
g23691(1) = AND(g14731, g20993)
g22316(1) = AND(g2837, g20270)
g26122(1) = AND(g24557, g19762)
g24854(1) = OR(g21453, g24002)
g22145(1) = AND(g14555, g18832)
g26153(1) = AND(g24565, g19780)
g24420(1) = AND(g23997, g18980)
g26635(1) = AND(g25321, g20617)
g24879(1) = OR(g21465, g24009)
g25530(1) = AND(g23750, g21414)
g26711(1) = AND(g25446, g20713)
g25122(1) = AND(g23374, g20592)
g24645(1) = AND(g22639, g19709)
g26303(1) = AND(g2685, g25439)
g24698(1) = AND(g22664, g19761)
g24514(1) = NOR(g23619, g23657)
g26091(1) = AND(g1691, g25082)
g25108(1) = AND(g23345, g20576)
g23404(1) = AND(g20063, g20247)
g25982(1) = AND(g2351, g25008)
g26649(1) = NOR(g9037, g24732)
g27238(1) = OR(g25879, g24464)
g26252(1) = AND(g2283, g25309)
g24931(1) = AND(g23153, g20178)
g23387(1) = AND(g16506, g20211)
g23646(1) = AND(g16959, g20737)
g27182(1) = OR(g25818, g24410)
g24546(1) = AND(g22447, g19523)
g25937(1) = OR(g24406, g22216)
g25949(1) = AND(g24701, g19559)
g25536(1) = AND(g23770, g21431)
g27509(1) = OR(g26023, g24640)
g25904(1) = AND(g14001, g24791)
g26205(1) = AND(g2098, g25492)
g26311(1) = AND(g2527, g25400)
g24658(1) = AND(g22645, g19732)
g26051(1) = AND(g24896, g14169)
g27663(1) = OR(g26323, g24820)
g22752(1) = AND(g15792, g19612)
g23386(1) = AND(g20034, g20207)
g24503(1) = AND(g22225, g19409)
g25835(1) = OR(g25367, g23855)
g22489(1) = AND(g12954, g19386)
g23857(1) = AND(g19626, g7908)
g22525(1) = AND(g13006, g19411)
g27269(1) = AND(g25943, g19734)
g23690(1) = AND(g14726, g20978)
g27268(1) = AND(g25942, g19733)
g25152(1) = AND(g23383, g20626)
g26302(1) = AND(g2393, g25349)
g26361(1) = OR(g24674, g22991)
g22686(1) = AND(g19335, g19577)
g23775(1) = AND(g14872, g21267)
g25928(1) = AND(g25022, g23436)
g25113(1) = AND(g23346, g20577)
g26249(1) = AND(g1858, g25300)
g24923(1) = AND(g23129, g20167)
g26204(1) = AND(g1720, g25275)
g24497(1) = NOR(g23533, g23553)
g26778(1) = AND(g25501, g20923)
g24148(1) = NOR(g19268, g19338)
I22298(1) = OR(g20371, g20161, g20151)
g24609(8) = NAND(g22850, g22650)
g23825(2) = OR(g20705, g20781)
g22400(4) = NOR(g19345, g15718)
g22450(4) = NOR(g19345, g15724)
I22830(1) = OR(g21429, g21338, g21307)
g22585(2) = OR(g20915, g21061)
g24591(8) = NAND(g22833, g22642)
g25575(1) = OR(g24139, g24140)
I23163(1) = OR(g20982, g21127, g21193, g21256)
I22280(1) = OR(g20271, g20150, g20134)
I22912(1) = OR(g21555, g21364, g21357)
I23162(1) = OR(g19919, g19968, g20014, g20841)
g25577(1) = OR(g24143, g24144)
g25576(1) = OR(g24141, g24142)
I22267(1) = OR(g20236, g20133, g20111)
g22531(2) = OR(g20773, g20922)
I22852(1) = OR(g21459, g21350, g21339)
g24145(1) = NOR(g19402, g19422)
I22880(1) = OR(g21509, g21356, g21351)
I22958(1) = OR(g21603, g21386, g21365)
I26523(1) = OR(g20720, g20857, g20998, g21143)
I22760(2) = NAND(g11939, g21434)
g22984(1) = NAND(g20114, g2868)
g22853(1) = NAND(g20219, g2922)
g22836(1) = NAND(g18918, g2852)
I22683(2) = NAND(g11893, g21434)
I20222(1) = NAND(g16272, I20221)
I23119(1) = NAND(g20076, I23118)
g22874(1) = NAND(g18918, g2844)
g22712(1) = NAND(g18957, g2864)
g23010(1) = NAND(g20516, g2984)
g22941(1) = NAND(g20219, g2970)
I22972(2) = NAND(g9657, g19638)
g22852(1) = NAND(g18957, g2856)
I22944(2) = NAND(g9492, g19620)
g23195(1) = NAND(g20136, g37)
g22921(1) = NAND(g20219, g2950)
I22753(2) = NAND(g11937, g21434)
I22792(2) = NAND(g11956, g21434)
I22844(2) = NAND(g12113, g21228)
I22899(2) = NAND(g12193, g21228)
I20205(1) = NAND(g11147, I20203)
I22717(2) = NAND(g11916, g21434)
g23266(1) = NAND(g18918, g2894)
I22871(2) = NAND(g12150, g21228)
g22940(1) = NAND(g18918, g2860)
I20204(1) = NAND(g16246, I20203)
g23956(1) = NOR(g18957, g18918, g20136, g20114)
I22822(2) = NAND(g11978, g21434)
I22929(2) = NAND(g12223, g21228)
I20166(1) = NAND(g16246, I20165)
I20167(1) = NAND(g990, I20165)
g22755(1) = NAND(g20136, g18984)
g22668(1) = NAND(g20219, g2912)
g22875(1) = NAND(g20516, g2980)
I22892(2) = NAND(g12189, g21228)
I22799(2) = NAND(g11960, g21434)
g22754(1) = NAND(g20114, g19376)
I22864(2) = NAND(g12146, g21228)
g22902(1) = NAND(g18957, g2848)
g22661(1) = NAND(g20136, g94)
g22715(1) = NAND(g20114, g2999)
I23120(1) = NAND(g417, I23118)
I22965(2) = NAND(g12288, g21228)
I20188(1) = NAND(g16272, I20187)
I20189(1) = NAND(g1333, I20187)
I22936(2) = NAND(g12226, g21228)
g14677(2) = NAND(I16779, I16780)
g23281(1) = NAND(g18957, g2898)
g22839(1) = NAND(g20114, g2988)
I21976(2) = NAND(g7680, g19620)
g22688(1) = NAND(g20219, g2936)
g22838(1) = NAND(g20219, g2960)
I21992(2) = NAND(g7670, g19638)
g22666(1) = NAND(g18957, g2878)
I22710(2) = NAND(g11915, g21434)
g22651(1) = NAND(g20114, g2873)
g22638(1) = NAND(g18957, g2886)
g22405(1) = NOR(g18957, g20136, g20114)
g23210(1) = NAND(g18957, g2882)
g22713(1) = NAND(g20114, g2890)
g22757(1) = NAND(g20114, g7891)
g22837(1) = NAND(g20219, g2907)
I20223(1) = NAND(g11170, I20221)
g22643(1) = NAND(g20136, g18954)
g18881(1) = NOT(I19671)
g20049(1) = NOT(I20318)
g20557(1) = NOT(I20647)
g20652(1) = NOT(I20744)
g20654(1) = NOT(I20750)
g20763(1) = NOT(I20816)
g20899(1) = NOT(I20861)
g20901(1) = NOT(I20867)
g21176(1) = NOT(I20954)
g21245(1) = NOT(I20982)
g21270(1) = NOT(I20999)
g21292(1) = NOT(I21033)
g21698(1) = NOT(g18562)
g21727(1) = NOT(I21300)
g26875(1) = OR(g21652, g25575)
g26876(1) = OR(g21655, g25576)
g26877(1) = OR(g21658, g25577)
g24276(1) = OR(g23083, g18646)
g25604(1) = OR(g24717, g18115)
g25607(1) = OR(g24773, g18118)
g25736(1) = OR(g25536, g18785)
g24216(1) = OR(g23416, g18197)
g24232(1) = OR(g22686, g18228)
g25668(1) = OR(g24646, g18623)
g24344(1) = OR(g22145, g18787)
g24274(1) = OR(g23187, g18631)
g24340(1) = OR(g24016, g18770)
g25633(1) = OR(g24420, g18282)
g24259(1) = OR(g23008, g18312)
g25684(1) = OR(g24983, g18643)
g25613(1) = OR(g25181, g18140)
g24244(1) = OR(g23349, g18255)
g25621(1) = OR(g24523, g18205)
g24235(1) = OR(g22632, g18238)
g25619(1) = OR(g24961, g18193)
g25656(1) = OR(g24945, g18609)
g24236(1) = OR(g22489, g18241)
g26917(1) = OR(g26122, g18233)
g24337(1) = OR(g23540, g18754)
g24336(1) = OR(g24012, g18753)
g24250(1) = OR(g22633, g18295)
g24251(1) = OR(g22637, g18296)
g24239(1) = OR(g22752, g18250)
g26897(1) = OR(g26611, g18176)
g24353(1) = OR(g23682, g18822)
g21903(1) = NOT(I21480)
g24253(1) = OR(g22525, g18300)
g24281(1) = OR(g23397, g18656)
g24237(1) = OR(g22515, g18242)
g25655(1) = OR(g24645, g18607)
g24269(1) = OR(g23131, g18613)
g28090(1) = OR(g27275, g18733)
g24209(1) = OR(g23415, g18122)
g24206(1) = OR(g23386, g18110)
g25669(1) = OR(g24657, g18624)
g24350(1) = OR(g23755, g18806)
g24210(1) = OR(g22900, g18125)
g28084(1) = OR(g27254, g18698)
g25625(1) = OR(g24553, g18226)
g25748(1) = OR(g25078, g18799)
g26899(1) = OR(g26844, g18199)
g25622(1) = OR(g24546, g18217)
g25749(1) = OR(g25094, g18800)
g25601(1) = OR(g24660, g18112)
g26915(1) = OR(g25900, g18230)
g25750(1) = OR(g25543, g18802)
g25721(1) = OR(g25057, g18766)
g24205(1) = OR(g23006, g18109)
g25763(1) = OR(g25113, g18817)
g24242(1) = OR(g22834, g18253)
g24245(1) = OR(g22849, g18256)
g24278(1) = OR(g23201, g18648)
g24282(1) = OR(g23407, g18657)
g26894(1) = OR(g25979, g18129)
g25654(1) = OR(g24634, g18606)
g25629(1) = OR(g24962, g18258)
g24262(1) = OR(g23387, g18315)
g25720(1) = OR(g25042, g18765)
g24261(1) = OR(g22862, g18314)
g25747(1) = OR(g25130, g18795)
g26922(1) = OR(g25902, g18288)
g25627(1) = OR(g24503, g18247)
g24254(1) = OR(g23265, g18306)
g24277(1) = OR(g23188, g18647)
g25603(1) = OR(g24698, g18114)
g25608(1) = OR(g24643, g18120)
g25611(1) = OR(g24931, g18128)
g26932(1) = OR(g26684, g18549)
g25624(1) = OR(g24408, g18224)
g21902(1) = NOT(I21477)
g28045(1) = OR(g27378, g18141)
g24208(1) = OR(g23404, g18121)
g24213(1) = OR(g23220, g18186)
g26898(1) = OR(g26387, g18194)
g25618(1) = OR(g25491, g18192)
g25600(1) = OR(g24650, g18111)
g26933(1) = OR(g26808, g18551)
g24268(1) = OR(g23025, g18612)
g24203(1) = OR(g22982, g18107)
g24346(1) = OR(g23725, g18789)
g24207(1) = OR(g23396, g18119)
g24348(1) = OR(g22149, g18804)
g28089(1) = OR(g27269, g18731)
g24233(1) = OR(g22590, g18236)
g25667(1) = OR(g24682, g18619)
g25612(1) = OR(g24941, g18132)
g26923(1) = OR(g25923, g18290)
g24211(1) = OR(g23572, g18138)
g24341(1) = OR(g23564, g18771)
g24201(1) = OR(g22848, g18104)
g24243(1) = OR(g22992, g18254)
g24335(1) = OR(g22165, g18678)
g25610(1) = OR(g24923, g18127)
g25606(1) = OR(g24761, g18117)
g28085(1) = OR(g27263, g18700)
g25722(1) = OR(g25530, g18768)
g25605(1) = OR(g24743, g18116)
g24272(1) = OR(g23056, g18629)
g24214(1) = OR(g23471, g18195)
g24355(1) = OR(g23799, g18824)
g24238(1) = OR(g23254, g18248)
g26895(1) = OR(g26783, g18148)
g24347(1) = OR(g23754, g18790)
g26921(1) = OR(g25955, g18285)
g28083(1) = OR(g27249, g18689)
g24212(1) = OR(g23280, g18155)
g25761(1) = OR(g25152, g18812)
g26931(1) = OR(g26778, g18547)
g26924(1) = OR(g26153, g18291)
g28087(1) = OR(g27255, g18720)
g25609(1) = OR(g24915, g18126)
g21722(1) = NOT(I21285)
g26930(1) = OR(g26799, g18544)
g24267(1) = OR(g23439, g18611)
g24249(1) = OR(g22624, g18294)
g28086(1) = OR(g27268, g18702)
g24270(1) = OR(g23165, g18614)
g25615(1) = OR(g24803, g18162)
g25617(1) = OR(g25466, g18189)
g24247(1) = OR(g22623, g18259)
g24215(1) = OR(g23484, g18196)
g25719(1) = OR(g25089, g18761)
g24231(1) = OR(g22589, g18201)
g25639(1) = OR(g25122, g18530)
g25614(1) = OR(g24797, g18161)
g24279(1) = OR(g23218, g15105)
g25708(1) = OR(g25526, g18751)
g24334(1) = OR(g23991, g18676)
g26929(1) = OR(g26635, g18543)
g24263(1) = OR(g23497, g18529)
g26912(1) = OR(g25946, g18209)
g24204(1) = OR(g22990, g18108)
g21723(1) = NOT(I21288)
g24275(1) = OR(g23474, g18645)
g24349(1) = OR(g23646, g18805)
g25634(1) = OR(g24559, g18284)
g25630(1) = OR(g24532, g18263)
g26927(1) = OR(g26711, g18539)
g25631(1) = OR(g24554, g18275)
g26896(1) = OR(g26341, g18171)
g25602(1) = OR(g24673, g18113)
g26916(1) = OR(g25916, g18232)
g24200(1) = OR(g22831, g18103)
g25764(1) = OR(g25551, g18819)
g24246(1) = OR(g23372, g18257)
g24255(1) = OR(g22835, g18308)
g24248(1) = OR(g22710, g18286)
g24234(1) = OR(g22622, g18237)
g25628(1) = OR(g24600, g18249)
g26934(1) = OR(g26845, g18556)
g24202(1) = OR(g22899, g18106)
g26919(1) = OR(g25951, g18267)
g24354(1) = OR(g23775, g18823)
g25636(1) = OR(g24507, g18305)
g26914(1) = OR(g25949, g18227)
g25670(1) = OR(g24967, g18626)
g25626(1) = OR(g24499, g18235)
g25762(1) = OR(g25095, g18816)
g24352(1) = OR(g22157, g18821)
g24342(1) = OR(g23691, g18772)
g21905(1) = NOT(I21486)
g24351(1) = OR(g23774, g18807)
g25637(1) = OR(g24618, g18307)
g25735(1) = OR(g25077, g18783)
g28088(1) = OR(g27264, g18729)
g24273(1) = OR(g23166, g18630)
g26928(1) = OR(g26713, g18541)
g25683(1) = OR(g24669, g18641)
g24258(1) = OR(g22851, g18311)
g25707(1) = OR(g25041, g18749)
g24339(1) = OR(g23690, g18756)
g21724(1) = NOT(I21291)
g25733(1) = OR(g25108, g18778)
g25638(1) = OR(g24977, g18316)
g24345(1) = OR(g23606, g18788)
g25635(1) = OR(g24504, g18293)
g25734(1) = OR(g25058, g18782)
g25653(1) = OR(g24664, g18602)
g21725(1) = NOT(I21294)
g25681(1) = OR(g24710, g18636)
g25705(1) = OR(g25069, g18744)
g24260(1) = OR(g23373, g18313)
g21726(1) = NOT(I21297)
g25682(1) = OR(g24658, g18640)
g25706(1) = OR(g25030, g18748)
g24338(1) = OR(g23658, g18755)
g21904(1) = NOT(I21483)
g24343(1) = OR(g23724, g18773)
g24252(1) = OR(g22518, g18299)
g24271(1) = OR(g23451, g18628)
g23499(1) = NOT(g20785)
g22494(1) = NOT(g19801)
g23611(1) = NOT(g18833)
g23988(1) = NOT(g19277)
g23924(1) = NOT(g18997)
g22182(7) = NOT(I21766)
g23432(1) = NOT(g21514)
g21271(1) = NOT(I21002)
g23271(1) = NOT(g20785)
g22155(1) = NOT(g19074)
g22170(1) = NOT(g19210)
g23461(1) = NOT(g18833)
g23031(1) = NOT(g19801)
g20653(1) = NOT(I20747)
g23887(1) = NOT(g18997)
g22167(1) = NOT(g19074)
g22194(2) = NOT(I21776)
g20558(1) = NOT(I20650)
g23528(1) = NOT(g18833)
g23843(1) = NOT(g19147)
g23869(1) = NOT(g19277)
g22763(66) = NOT(I22046)
g28294(1) = NOT(g27295)
g23868(1) = NOT(g19277)
g20655(1) = NOT(I20753)
g24156(1) = NOT(I23312)
g23259(1) = NOT(g21070)
g22305(1) = NOT(g19801)
g23258(1) = NOT(g20924)
g23244(1) = NOT(I22343)
g22177(1) = NOT(g19074)
g19862(2) = NOT(I20233)
g23375(1) = NOT(g20924)
g24264(1) = OR(g22310, g18559)
g23879(1) = NOT(g19210)
g23970(1) = NOT(g19277)
g23878(1) = NOT(g19147)
g23337(1) = NOT(g20924)
g23886(1) = NOT(g21468)
g22166(1) = NOT(g18997)
g23792(1) = NOT(g19074)
g23967(1) = NOT(g19210)
g23994(1) = NOT(g19277)
g23459(1) = NOT(g21611)
g23458(1) = NOT(I22583)
g22907(1) = NOT(g20453)
g23545(1) = NOT(g21562)
g23444(1) = NOT(I22561)
I21934(1) = NOT(g21273)
g23086(1) = NOT(g20283)
g27014(1) = NOT(g25888)
g23322(1) = NOT(I22425)
g22519(1) = NOT(g19801)
g22176(1) = NOT(g18997)
g25228(1) = NOT(g23828)
g22154(1) = NOT(g19074)
g22935(1) = NOT(g20283)
g23353(1) = NOT(g20924)
g22883(1) = NOT(g20391)
I22989(1) = NOT(g21175)
g23336(1) = NOT(g20924)
g23966(1) = NOT(g19210)
g22215(1) = NOT(g19277)
g23017(1) = NOT(g20453)
g23289(1) = NOT(g20924)
g24373(1) = NOT(g22908)
g22906(1) = NOT(g20453)
g22546(1) = NOT(I21918)
g23571(1) = NOT(g18833)
g23495(1) = NOT(I22622)
g23985(1) = NOT(g19210)
I22788(1) = NOT(g18940)
g24000(1) = NOT(g19277)
g23260(1) = NOT(g21070)
g23842(1) = NOT(g19147)
g23384(1) = NOT(I22485)
g23489(1) = NOT(g21468)
g24568(1) = NOT(g22942)
g23559(1) = NOT(g21070)
g23525(1) = NOT(g21562)
g23488(1) = NOT(g21468)
g23016(1) = NOT(g20453)
g23558(1) = NOT(g20924)
g22200(1) = NOT(g19277)
g23893(1) = NOT(g19074)
g23544(1) = NOT(g21562)
g22683(1) = NOT(I22000)
g23610(1) = NOT(g18833)
g22973(1) = NOT(g20330)
g23270(1) = NOT(g20785)
g23460(1) = NOT(g21611)
g23939(1) = NOT(g19074)
g23030(1) = NOT(g20453)
g23938(1) = NOT(g18997)
g23875(1) = NOT(g18997)
g25080(1) = NOT(g23742)
g23219(1) = NOT(I22316)
g22214(1) = NOT(g19210)
g22207(1) = NOT(I21787)
g23915(1) = NOT(g19277)
g23277(1) = NOT(I22380)
g23494(1) = NOT(I22619)
g24818(1) = NOT(g23191)
g23984(1) = NOT(g19210)
g23419(1) = NOT(g21468)
g23352(1) = NOT(g20924)
g25225(1) = NOT(g23802)
g22882(1) = NOT(g20391)
g28608(1) = NOT(g27670)
g23418(1) = NOT(g21468)
g27492(1) = NOT(g26598)
g25244(1) = NOT(g23802)
g23589(1) = NOT(g21468)
g23524(1) = NOT(g21562)
g23477(1) = NOT(g21468)
g22758(1) = NOT(g20330)
g24372(1) = NOT(g22885)
g23864(1) = NOT(g19210)
g23022(1) = NOT(g20283)
g23749(1) = NOT(g18997)
g23313(1) = NOT(g21070)
g25994(1) = NOT(g24575)
g24516(1) = NOT(g22670)
g23305(1) = NOT(g20391)
g29172(1) = NOT(g27020)
g24266(1) = OR(g22329, g18561)
g21177(1) = NOT(I20957)
g22332(5) = NOT(I21838)
I22785(1) = NOT(g18940)
g23874(1) = NOT(g18997)
g23665(1) = NOT(g21562)
g23320(1) = NOT(I22419)
g23450(1) = NOT(I22571)
g23476(1) = NOT(g21468)
g23485(1) = NOT(g20785)
g23555(2) = NOT(I22692)
g23570(1) = NOT(g18833)
g23914(1) = NOT(g19210)
g24153(1) = NOT(I23303)
g23907(1) = NOT(g19074)
g23567(1) = NOT(g21562)
g23238(1) = NOT(g20924)
g28441(1) = NOT(g27629)
g23941(1) = NOT(g19074)
g23519(1) = NOT(g21468)
g23518(1) = NOT(g21070)
g23154(7) = NOT(I22264)
g23935(1) = NOT(g19210)
g22976(2) = NOT(I22149)
g22923(2) = NOT(I22124)
g22541(1) = NOT(I21911)
g23215(1) = NOT(g20785)
g23501(1) = NOT(g20924)
g22358(1) = NOT(g19801)
g23906(1) = NOT(g19074)
g23284(1) = NOT(g20785)
g23304(1) = NOT(g20785)
g23566(1) = NOT(g21562)
g22173(2) = NOT(I21757)
g24522(1) = NOT(g22689)
g27046(3) = NOR(g7544, g25888)
g23138(1) = NOT(g20453)
g23333(1) = NOT(g20785)
I22889(1) = NOT(g18926)
g23963(1) = NOT(g19147)
g22927(1) = NOT(I22128)
g22409(8) = NOT(I21860)
g23585(1) = NOT(g21070)
g23609(1) = NOT(g21611)
g24397(1) = NOT(g22908)
g22903(1) = NOT(g20330)
g23312(1) = NOT(g21070)
g23608(1) = NOT(g21611)
g24509(1) = NOT(g22689)
I26296(1) = NOT(g26820)
g22981(1) = NOT(g20283)
g20900(1) = NOT(I20864)
g23813(1) = NOT(g18997)
g27463(3) = NAND(g287, g26330, g23204)
g22898(1) = NOT(g20283)
g23732(1) = NOT(g18833)
g23013(1) = NOT(g20330)
g23214(1) = NOT(g20785)
g22926(1) = NOT(g20391)
g23539(1) = NOT(g21070)
g23005(1) = NOT(g20283)
g23538(1) = NOT(g20924)
g24152(1) = NOT(I23300)
g24396(1) = NOT(g22885)
g22997(1) = NOT(g20391)
g27059(3) = NOR(g7577, g25895)
g23235(1) = NOT(g20785)
g22360(9) = NOT(I21849)
g28648(1) = NOT(g27693)
g23515(1) = NOT(g20785)
g23882(1) = NOT(g19277)
g23414(1) = NOT(I22525)
g22220(2) = NOT(I21802)
g28633(1) = NOT(g27687)
I22886(1) = NOT(g18926)
g22147(1) = NOT(g18997)
g23435(1) = NOT(g18833)
g23360(1) = NOT(I22461)
g22151(1) = NOT(I21734)
g23849(1) = NOT(g19277)
g22996(1) = NOT(g20330)
g23940(1) = NOT(g19074)
g23399(1) = NOT(g21514)
g23848(1) = NOT(g19210)
g23398(1) = NOT(g21468)
g24003(1) = NOT(g21514)
g23263(1) = NOT(I22366)
g22319(5) = NOT(I21831)
g23332(1) = NOT(g20785)
g22227(1) = NOT(g19801)
g23406(1) = NOT(g20330)
g23962(1) = NOT(g19147)
g23361(1) = NOT(I22464)
g23500(1) = NOT(g20924)
g23004(1) = NOT(g20283)
g23221(1) = NOT(g20785)
g22957(15) = NOT(I22143)
I22748(1) = NOT(g19458)
g22146(1) = NOT(g18997)
g23947(1) = NOT(g19210)
g23273(1) = NOT(g21070)
g22698(8) = NOT(I22009)
g23812(1) = NOT(g18997)
g24505(1) = NOT(g22689)
g24404(1) = NOT(g22908)
g23507(1) = NOT(g21562)
g27528(3) = NOR(g8770, g26352, g11083)
I22180(1) = NOT(g21366)
g23421(1) = NOT(g21562)
g23012(1) = NOT(g20330)
g23541(1) = NOT(g21514)
g23473(1) = NOT(g20785)
g23788(1) = NOT(g18997)
g23359(1) = NOT(I22458)
g23321(1) = NOT(I22422)
g22980(1) = NOT(I22153)
I22557(1) = NOT(g20695)
g23434(1) = NOT(g21611)
g23946(1) = NOT(g19210)
g22181(1) = NOT(g19277)
g28144(2) = AND(g4608, g27020)
g23291(1) = NOT(g21070)
g22520(1) = NOT(g19801)
g20050(1) = NOT(I20321)
g23029(1) = NOT(g20453)
g23506(1) = NOT(g21514)
g23028(1) = NOT(g20391)
g23202(1) = NOT(I22302)
g22987(1) = NOT(g20391)
g23927(1) = NOT(g19074)
g22658(1) = NOT(I21969)
g23649(1) = NOT(g18833)
g22339(1) = NOT(g19801)
g23648(1) = NOT(g18833)
g22338(1) = NOT(g19801)
g23491(1) = NOT(g21514)
g23903(1) = NOT(g18997)
g25013(1) = NOT(g23599)
g24548(1) = NOT(g22942)
g22197(1) = NOT(g19074)
g22855(1) = NOT(g20391)
g23767(1) = NOT(g18997)
g23794(1) = NOT(g19147)
g23395(1) = NOT(I22502)
g23899(1) = NOT(g19277)
g22867(1) = NOT(g20391)
g23898(1) = NOT(g19277)
g24533(1) = NOT(g22876)
g23521(1) = NOT(g21468)
g23232(1) = NOT(I22331)
g22202(5) = NOT(I21784)
g22979(1) = NOT(g20453)
g23861(1) = NOT(g19147)
g23247(1) = NOT(g20924)
g22986(1) = NOT(g20330)
g25026(1) = AND(g22929, g10503)
g23926(1) = NOT(g19074)
I22745(1) = NOT(g19458)
g23388(1) = NOT(g21070)
g23534(2) = NOT(I22665)
g23272(1) = NOT(g20924)
g23462(8) = NOT(I22589)
g23032(8) = NOT(I22211)
g22526(1) = NOT(g19801)
g23061(1) = NOT(g20283)
g22866(1) = NOT(g20330)
g23447(1) = NOT(g21562)
g23362(1) = NOT(I22467)
g23629(1) = NOT(g21514)
g22300(2) = NOT(I21815)
g27017(1) = NOT(g25895)
g21246(1) = NOT(I20985)
g23246(1) = NOT(g20785)
g20764(1) = NOT(I20819)
g23355(1) = NOT(g21070)
g23859(1) = NOT(g19074)
g22854(1) = NOT(g20330)
g23858(1) = NOT(g18997)
g23172(9) = NOT(I22275)
g23394(1) = NOT(I22499)
g22456(1) = NOT(g19801)
g23420(1) = NOT(g21514)
I21922(1) = NOT(g21335)
g23446(1) = NOT(g21562)
g23227(1) = NOT(g20924)
g23059(1) = NOT(g20453)
g22721(1) = NOT(I22028)
g23058(1) = NOT(g20453)
g22341(1) = NOT(g19801)
g22156(1) = NOT(g19147)
g23902(1) = NOT(g21468)
g23301(1) = NOT(g21037)
g23377(1) = NOT(g21070)
g22180(1) = NOT(g19210)
g24010(1) = NOT(g21562)
g23290(1) = NOT(g20924)
g23698(1) = NOT(g21611)
g23427(1) = NOT(I22542)
g22210(2) = NOT(I21792)
g24159(1) = NOT(I23321)
g23403(1) = NOT(I22512)
g23547(1) = NOT(g21611)
g23895(1) = NOT(g19147)
g24158(1) = NOT(I23318)
g23226(1) = NOT(g20924)
g23481(1) = NOT(I22604)
g22975(1) = NOT(g20391)
g23252(1) = NOT(I22353)
g23490(1) = NOT(g21514)
g24017(1) = NOT(g18833)
g23376(1) = NOT(g21070)
g23385(1) = NOT(I22488)
g23354(1) = NOT(g20453)
g22169(1) = NOT(g19147)
g22884(1) = NOT(g20453)
g23888(1) = NOT(g18997)
g28307(1) = NOT(g27306)
g22168(1) = NOT(g19147)
I26925(1) = NOT(g27015)
g24571(1) = NOT(g22942)
g25423(1) = NOT(I24558)
g23426(1) = NOT(I22539)
g23520(1) = NOT(g21468)
g22223(1) = NOT(g19210)
g23546(1) = NOT(g21611)
g23088(14) = NOT(I22240)
g22922(1) = NOT(g20330)
g23860(1) = NOT(g19074)
g22179(1) = NOT(g19210)
g24997(1) = AND(g22929, g10419)
g22178(1) = NOT(g19147)
g23987(1) = NOT(g19277)
g23250(1) = NOT(g21070)
g24525(1) = NOT(g22670)
g22936(1) = NOT(g20283)
g23339(1) = NOT(g21070)
g23943(1) = NOT(g19147)
g23338(1) = NOT(g20453)
g23969(1) = NOT(g19277)
g23968(1) = NOT(g18833)
g21293(1) = NOT(I21036)
g23527(1) = NOT(g21611)
g22543(1) = NOT(g19801)
g23503(1) = NOT(g21468)
g23894(1) = NOT(g19074)
g25032(1) = NOT(g23639)
g23819(1) = NOT(g19147)
g27654(3) = NAND(g164, g26598, g23042)
g23257(1) = NOT(g20924)
g23111(1) = NOT(g20391)
g22974(1) = NOT(g20330)
g23986(1) = NOT(g18833)
g24160(1) = NOT(I23324)
g22841(1) = NOT(g20391)
g23877(1) = NOT(g19147)
g28321(1) = NOT(g27317)
g25246(1) = NOT(g23828)
g23196(1) = NOT(g20785)
g23018(1) = NOT(g19801)
g23526(1) = NOT(g21611)
g24623(1) = NOT(g23076)
g23457(1) = NOT(I22580)
g24155(1) = NOT(I23309)
g22493(1) = NOT(g19801)
g23001(1) = NOT(g19801)
g23256(1) = NOT(g20785)
g23923(1) = NOT(g18997)
g23300(1) = NOT(g20283)
g24524(1) = NOT(g22876)
g27349(1) = NOT(g26352)
g23066(1) = NOT(g20330)
g23876(1) = NOT(g19074)
g25044(1) = NOT(g23675)
g23511(1) = NOT(I22640)
g23230(1) = NOT(I22327)
g23456(1) = NOT(g21514)
g24560(1) = NOT(g22942)
g23480(1) = NOT(I22601)
g23916(1) = NOT(g19277)
g23307(1) = NOT(g20924)
g23243(1) = NOT(g21070)
g23431(1) = NOT(g21514)
g26081(1) = NOT(g24619)
g23942(1) = NOT(g21562)
g23335(1) = NOT(g20391)
g23839(1) = NOT(g18997)
g23930(1) = NOT(g19147)
g23993(1) = NOT(g19277)
g23838(1) = NOT(g18997)
g23965(1) = NOT(g21611)
g22542(1) = NOT(g19801)
g23487(1) = NOT(g20924)
g23502(1) = NOT(g21070)
g23443(1) = NOT(g21468)
g23279(1) = NOT(g21037)
g22905(1) = NOT(I22114)
g24154(1) = NOT(I23306)
g23278(1) = NOT(g20283)
g22593(1) = NOT(g19801)
g23306(1) = NOT(g20924)
g23815(1) = NOT(g19074)
g22153(1) = NOT(g18997)
g22635(1) = NOT(g19801)
g23937(1) = NOT(g19277)
g23410(1) = NOT(g21562)
g23479(1) = NOT(g21562)
g23363(8) = NOT(I22470)
g23478(1) = NOT(g21514)
g23015(1) = NOT(g20391)
I25530(1) = NOT(g25222)
g23486(1) = NOT(g20785)
I26638(1) = NOT(g27965)
g25060(1) = NOT(g23708)
g25197(1) = NOT(g23958)
g22303(1) = NOT(g19277)
g24636(1) = NOT(g23121)
g23922(1) = NOT(g18997)
g23953(1) = NOT(g19277)
g22840(1) = NOT(g20330)
g23417(1) = NOT(g20391)
g23936(1) = NOT(g19210)
g22647(1) = NOT(I21959)
g22192(1) = NOT(g19801)
g23334(1) = NOT(g20785)
g23964(1) = NOT(g19147)
g23216(1) = NOT(g20924)
g23543(1) = NOT(g21514)
g22904(1) = NOT(I22111)
g23000(1) = NOT(g20453)
g23569(1) = NOT(g21611)
g23568(1) = NOT(g21611)
g23242(1) = NOT(g21070)
g22847(1) = NOT(g20283)
g23814(1) = NOT(g19074)
g24013(1) = NOT(g21611)
g18882(1) = NOT(I19674)
g23841(1) = NOT(g19074)
g23992(1) = NOT(g19210)
g23510(1) = NOT(g18833)
g22213(1) = NOT(g19147)
g23014(1) = NOT(g20391)
g22592(1) = NOT(I21930)
g24515(1) = NOT(g22689)
g23430(1) = NOT(I22547)
g20902(1) = NOT(I20870)
g23493(1) = NOT(g21611)
g23237(1) = NOT(g20924)
g23340(1) = NOT(g21070)
g23983(1) = NOT(g19210)
g23517(1) = NOT(g21070)
g22928(1) = NOT(I22131)
g23523(1) = NOT(g21514)
g23863(1) = NOT(g19210)
g23222(1) = NOT(g20785)
g23347(1) = NOT(I22444)
g23253(1) = NOT(g21037)
g24361(1) = NOT(g22885)
g25210(1) = NOT(g23802)
g23236(1) = NOT(g20785)
g23952(1) = NOT(g19277)
g23351(1) = NOT(g20924)
g22881(1) = NOT(I22096)
g23821(1) = NOT(g19210)
g23264(1) = NOT(g21037)
g23516(1) = NOT(g20924)
I22031(1) = NOT(g21387)
g23422(1) = NOT(g21611)
g23542(1) = NOT(g21514)
g23021(1) = NOT(g20283)
g23913(1) = NOT(g19147)
g22999(1) = NOT(g20453)
g23607(1) = NOT(g21611)
g23905(1) = NOT(g21514)
g23274(1) = NOT(g21070)
g22998(1) = NOT(g20391)
g23565(1) = NOT(g21562)
g23409(1) = NOT(g21514)
g23408(1) = NOT(g21468)
g24535(1) = NOT(g22942)
g22148(1) = NOT(g19074)
g23537(1) = NOT(g20785)
g23283(1) = NOT(g20785)
g23492(1) = NOT(g21562)
g23303(1) = NOT(g20785)
g24265(1) = OR(g22316, g18560)
g23982(1) = NOT(g19147)
g23840(1) = NOT(g19074)
g23390(1) = NOT(g21468)
I21810(1) = NOT(g20596)
g24648(1) = NOT(g23148)
g23522(1) = NOT(g21514)
g25230(1) = NOT(g23314)
g23483(1) = NOT(g18833)
g23862(1) = NOT(g19147)
g23904(1) = NOT(g18997)
g23847(1) = NOT(g19210)
g23509(1) = NOT(g21611)
g28620(1) = NOT(g27679)
g24389(1) = NOT(g22908)
g23508(1) = NOT(g21562)
g24388(1) = NOT(g22885)
g22317(1) = NOT(g19801)
g24534(1) = NOT(g22670)
g22626(5) = NOT(I21941)
g23452(1) = NOT(g21468)
g23912(1) = NOT(g19147)
g22856(1) = NOT(g20453)
g22995(1) = NOT(g20330)
g23350(1) = NOT(g20785)
g23820(1) = NOT(g19147)
g23152(1) = NOT(g20283)
g22989(1) = NOT(g20453)
g23929(1) = NOT(g19147)
g22988(1) = NOT(g20391)
g23928(1) = NOT(g21562)
g25264(1) = NOT(g23828)
g23046(1) = NOT(g20283)
g23787(1) = NOT(g18997)
g21282(1) = NOT(I21019)
g23282(1) = NOT(g20330)
g23302(1) = NOT(g20330)
g22199(1) = NOT(g19210)
g22198(1) = NOT(g19147)
g22528(1) = NOT(g19801)
g23769(1) = NOT(g19074)
g22330(1) = NOT(g19801)
g23768(1) = NOT(g18997)
g24540(1) = NOT(g22942)
g22868(1) = NOT(g20453)
g23881(1) = NOT(g19277)
g23027(1) = NOT(g20391)
g23299(1) = NOT(I22400)
g23249(1) = NOT(g21070)
g23482(1) = NOT(g18833)
g23248(1) = NOT(g20924)
g24374(1) = OR(g19345, g24004)
g23647(1) = NOT(g18833)
g23945(1) = NOT(g21611)
g23356(1) = NOT(g21070)
g23999(1) = NOT(g21468)
g23233(1) = NOT(g21037)
I22177(1) = NOT(g21366)
g23449(1) = NOT(g18833)
g23897(1) = NOT(g19210)
g23448(1) = NOT(g21611)
g23961(1) = NOT(g19074)
g23505(1) = NOT(g21514)
g24385(1) = NOT(g22908)
g23026(1) = NOT(g20391)
g27018(1) = NOT(I25750)
g22159(1) = NOT(I21744)
g23433(1) = NOT(g21562)
g22144(1) = NOT(g18997)
g27597(1) = NOT(g26745)
g23896(1) = NOT(g19210)
g22224(1) = NOT(g19277)
g23228(1) = NOT(g21070)
g23011(1) = NOT(g20330)
g22495(1) = NOT(g19801)
g23582(2) = NOT(I22729)
g22985(1) = NOT(g20330)
g23925(1) = NOT(g21514)
g23378(1) = NOT(g21070)
g24527(1) = NOT(g22670)
g23944(1) = NOT(g19147)
g25213(1) = NOT(g23293)
g27717(2) = NOR(g9492, g26745)
g23429(1) = NOT(g20453)
g23793(1) = NOT(g19074)
g22830(1) = NOT(g20283)
g23549(1) = NOT(g18833)
g22865(1) = NOT(g20330)
g23548(1) = NOT(g18833)
g23504(1) = NOT(g21468)
g24384(1) = NOT(g22885)
g28500(3) = NAND(g590, g27629, g12323)
g22189(1) = NOT(I21769)
g23057(1) = NOT(g20453)
g23128(1) = NOT(g20283)
g23245(1) = NOT(g20785)
g23323(1) = NOT(g20283)
g24526(1) = NOT(g22942)
g27277(1) = AND(g26359, g14191)
g27279(1) = NOT(g26330)
g23995(1) = NOT(g19277)
g23880(1) = NOT(g19210)
g22455(1) = NOT(g19801)
g28669(1) = NOT(g27705)
g22201(1) = NOT(g19277)
g23445(1) = NOT(I22564)
g24157(1) = NOT(I23315)
g22075(1) = AND(g6247, g19210)
g21989(1) = AND(g5587, g19074)
g26826(1) = AND(g24907, g15747)
g22037(1) = AND(g5941, g19147)
g27363(1) = AND(g10231, g26812)
g21988(1) = AND(g5583, g19074)
g21924(1) = AND(g5057, g21468)
g21753(1) = AND(g3179, g20785)
g25482(2) = AND(g5752, g23816, I24597)
I24684(1) = AND(g20014, g24033, g24034, g24035)
g21736(1) = AND(g3065, g20330)
g21887(1) = AND(g15101, g19801)
g27572(1) = OR(g26129, g24724)
g21843(1) = AND(g3869, g21070)
g21764(1) = AND(g3227, g20785)
I27528(1) = AND(g20998, g24118, g24119, g24120)
g28686(1) = AND(g27574, g20650)
g22119(1) = AND(g6581, g19277)
g21869(1) = AND(g4087, g19801)
g21960(1) = AND(g5421, g21514)
g27676(1) = AND(g26377, g20627)
g27685(1) = AND(g13032, g25895)
g22118(1) = AND(g6605, g19277)
g21868(1) = AND(g4076, g19801)
g22022(1) = AND(g5873, g19147)
g21709(1) = AND(g283, g20283)
g27334(1) = AND(g12539, g26769)
g28219(1) = AND(g9316, g27573)
g21708(1) = AND(g15049, g20283)
g22053(1) = AND(g6116, g21611)
g25956(1) = NOR(g1413, g24609)
g22036(1) = AND(g5937, g19147)
g22101(1) = AND(g6474, g18833)
g27289(1) = OR(g25925, g25927)
g21810(1) = AND(g3578, g20924)
g21774(1) = AND(g3361, g20391)
g28617(1) = AND(g27533, g20552)
g21955(1) = AND(g5385, g21514)
g22064(1) = AND(g15162, g19210)
g21879(1) = AND(g4132, g19801)
g21970(1) = AND(g5401, g21514)
g21878(1) = AND(g4129, g19801)
g22536(1) = NOR(g1379, g19720)
g21886(1) = AND(g4153, g19801)
g21792(1) = AND(g3396, g20391)
g22009(1) = AND(g5782, g21562)
g21967(1) = AND(g5456, g21514)
g21994(1) = AND(g5607, g19074)
g22008(1) = AND(g5774, g21562)
g28352(1) = AND(g10014, g27705)
g21919(1) = AND(g15144, g21468)
g27230(1) = AND(g25906, g19558)
g27293(1) = AND(g9972, g26655)
g21918(1) = AND(g5097, g21468)
g22074(1) = AND(g6239, g19210)
g21817(1) = AND(g3606, g20924)
g22545(1) = NOR(g1373, g19720)
g21977(1) = AND(g5535, g19074)
g22092(1) = AND(g6419, g18833)
g21783(1) = AND(g3419, g20391)
I27509(1) = AND(g24084, g24085, g24086, g24087)
g21823(1) = AND(g3731, g20453)
g27041(1) = AND(g8519, g26330)
g21966(1) = AND(g5406, g21514)
g27340(1) = AND(g10199, g26784)
g26348(1) = OR(g8466, g24609)
g27684(1) = AND(g26386, g20657)
g28642(1) = AND(g27555, g20598)
g22083(1) = AND(g6287, g19210)
g28630(1) = AND(g27544, g20575)
g26080(1) = OR(g19393, g24502)
g21816(1) = AND(g3602, g20924)
g21976(1) = AND(g5527, g19074)
g21985(1) = AND(g5571, g19074)
g28555(1) = AND(g27429, g20373)
g21752(1) = AND(g3171, g20785)
g28570(1) = AND(g27456, g20434)
g27590(1) = OR(g26179, g24764)
g21954(1) = AND(g5381, g21514)
g24908(2) = AND(g3752, g23239, I24075)
g28238(1) = AND(g27133, g19658)
g21842(1) = AND(g3863, g21070)
g27351(1) = AND(g10218, g26804)
g28154(1) = AND(g8492, g27306)
g21830(1) = AND(g3774, g20453)
g22399(1) = NOR(g1367, g19720)
g22115(1) = AND(g6573, g19277)
g21865(1) = AND(g3965, g21070)
g21713(1) = AND(g298, g20283)
g22052(1) = AND(g6113, g21611)
g21705(1) = AND(g209, g20283)
g28215(1) = AND(g9264, g27565)
g27208(1) = AND(g9037, g26598)
g21939(1) = AND(g5224, g18997)
g21938(1) = AND(g5216, g18997)
g28304(1) = AND(g27226, g19753)
g21875(1) = AND(g4116, g19801)
g22013(1) = AND(g5802, g21562)
g21837(1) = AND(g3719, g20453)
g26328(1) = OR(g1183, g24591)
g22005(1) = AND(g5759, g21562)
g27292(1) = AND(g1714, g26654)
g28333(1) = AND(g27239, g19787)
g21915(1) = AND(g5080, g21468)
g22100(1) = AND(g6466, g18833)
g21782(1) = AND(g3416, g20391)
g21984(1) = AND(g5563, g19074)
g28554(1) = AND(g27426, g20372)
g27327(1) = AND(g2116, g26732)
g21822(1) = AND(g3727, g20453)
g27303(1) = AND(g11996, g26681)
g21853(1) = AND(g3917, g21070)
g28813(1) = AND(g4104, g27038)
g21836(1) = AND(g3805, g20453)
g27569(1) = OR(g26124, g24721)
g22114(1) = AND(g6565, g19277)
g21864(1) = AND(g3961, g21070)
g22082(1) = AND(g6283, g19210)
g22107(1) = AND(g6411, g18833)
g21749(1) = AND(g3155, g20785)
g27578(1) = OR(g26155, g24747)
g21748(1) = AND(g15089, g20785)
g21704(1) = AND(g164, g20283)
g25459(2) = AND(g6058, g23844, I24582)
g21809(1) = AND(g3574, g20924)
g21808(1) = AND(g3570, g20924)
g27326(1) = AND(g12048, g26731)
g22135(1) = AND(g6657, g19277)
g21733(1) = AND(g3034, g20330)
g21874(1) = AND(g4112, g19801)
g25159(1) = AND(g4907, g22908)
g22049(1) = AND(g6082, g21611)
g25901(1) = AND(g24853, g16290)
g28235(1) = AND(g9467, g27592)
g22048(1) = AND(g6052, g21611)
I27514(1) = AND(g24091, g24092, g24093, g24094)
g22004(1) = AND(g5742, g21562)
g21712(1) = AND(g294, g20283)
g21914(1) = AND(g5077, g21468)
I24710(1) = AND(g24071, g24072, g24073, g24074)
g22106(1) = AND(g6497, g18833)
g21907(1) = AND(g5033, g21468)
g22033(1) = AND(g5925, g19147)
g21941(1) = AND(g5232, g18997)
g27311(1) = AND(g12431, g26693)
g27596(1) = OR(g26207, g24775)
I24694(1) = AND(g20982, g24047, g24048, g24049)
I24695(1) = AND(g24050, g24051, g24052, g24053)
g27970(1) = OR(g26514, g25050)
g21935(1) = AND(g5196, g18997)
g21883(1) = AND(g4141, g19801)
g22012(1) = AND(g5752, g21562)
I27504(1) = AND(g24077, g24078, g24079, g24080)
g27350(1) = AND(g10217, g26803)
g25374(2) = AND(g5366, g23789, I24527)
g21729(1) = AND(g3021, g20330)
g21728(1) = AND(g3010, g20330)
g19764(1) = NAND(I20166, I20167)
I27533(1) = AND(g21143, g24125, g24126, g24127)
g22121(1) = AND(g6593, g19277)
g21906(1) = AND(g5022, g21468)
g25488(2) = AND(g6404, g23865, I24603)
g25865(1) = AND(g25545, g18991)
g22134(1) = AND(g6653, g19277)
g22029(1) = AND(g5901, g19147)
g22028(1) = AND(g5893, g19147)
g27302(1) = AND(g1848, g26680)
g23796(3) = OR(g21462, g21433, I22958)
g21852(1) = AND(g3909, g21070)
g28812(1) = AND(g26972, g13037)
g25124(1) = AND(g4917, g22908)
g21963(1) = AND(g5436, g21514)
g25939(1) = AND(g24583, g19490)
g23198(3) = OR(g20214, g20199, I22298)
g21921(1) = AND(g5109, g21468)
g26822(1) = AND(g24841, g13116)
g22521(1) = NOR(g1036, g19699)
g21745(1) = AND(g3017, g20330)
g21799(1) = AND(g3530, g20924)
g21813(1) = AND(g3590, g20924)
g28541(1) = AND(g27403, g20274)
g27710(1) = AND(g26422, g20904)
g21798(1) = AND(g3522, g20924)
g21973(1) = AND(g5511, g19074)
g21805(1) = AND(g3550, g20924)
g25915(1) = AND(g24926, g9602)
g21732(1) = AND(g3004, g20330)
g21934(1) = AND(g5220, g18997)
g23687(3) = OR(g21384, g21363, I22830)
g21761(1) = AND(g3215, g20785)
I24690(1) = AND(g24043, g24044, g24045, g24046)
g26749(1) = AND(g24494, g23578)
g19792(1) = NAND(I20204, I20205)
g22448(1) = NOR(g1018, g19699)
g22045(1) = AND(g6069, g21611)
g22099(1) = AND(g6462, g18833)
g25944(1) = NOR(g7716, g24591)
g27331(1) = AND(g10177, g26754)
g22098(1) = AND(g6459, g18833)
g22032(1) = AND(g5921, g19147)
g21771(1) = AND(g3255, g20785)
g22061(1) = AND(g6065, g21611)
g23751(3) = OR(g21415, g21402, I22880)
g27723(1) = AND(g26512, g21049)
g21882(1) = AND(g4057, g19801)
g21991(1) = AND(g5595, g19074)
g27646(1) = AND(g13094, g25773)
g26712(1) = AND(g24508, g24463)
g22071(1) = AND(g6251, g19210)
g21759(1) = AND(g3199, g20785)
g21758(1) = AND(g3191, g20785)
g24881(2) = AND(g3050, g23211, I24048)
g21744(1) = AND(g3103, g20330)
g21849(1) = AND(g3889, g21070)
g21940(1) = AND(g5228, g18997)
g28247(1) = AND(g27147, g19675)
g21848(1) = AND(g3913, g21070)
g21804(1) = AND(g3542, g20924)
I24689(1) = AND(g20841, g24040, g24041, g24042)
g25948(1) = NOR(g7752, g24609)
g28612(1) = AND(g27524, g20539)
g28324(1) = AND(g9875, g27687)
g25950(1) = NOR(g1070, g24591)
g24799(3) = OR(g23901, g23921)
g24552(1) = AND(g22487, g19538)
I24674(1) = AND(g19919, g24019, g24020, g24021)
I24675(1) = AND(g24022, g24023, g24024, g24025)
g22059(1) = AND(g6148, g21611)
g21962(1) = AND(g5428, g21514)
g22025(1) = AND(g5905, g19147)
g22058(1) = AND(g6098, g21611)
g21833(1) = AND(g15096, g20453)
g24577(1) = OR(g2856, g22531)
g25518(2) = AND(g6444, g23865, I24625)
g22044(1) = AND(g6058, g21611)
I24709(1) = AND(g21256, g24068, g24069, g24070)
g22120(1) = AND(g6585, g19277)
g21947(1) = AND(g5256, g18997)
g24897(2) = AND(g3401, g23223, I24064)
g21812(1) = AND(g3586, g20924)
g27283(1) = OR(g25922, g25924)
g21951(1) = AND(g5272, g18997)
g21972(1) = AND(g15152, g19074)
g21795(1) = AND(g3506, g20924)
g28151(1) = AND(g8426, g27295)
g22127(1) = AND(g6625, g19277)
g24705(1) = OR(g2890, g23267)
g21789(1) = AND(g3451, g20391)
g21788(1) = AND(g3401, g20391)
g22103(1) = AND(g15164, g18833)
g21829(1) = AND(g3770, g20453)
g21920(1) = AND(g5062, g21468)
g22095(1) = AND(g6428, g18833)
g28318(1) = AND(g27233, g19770)
g28227(1) = AND(g9397, g27583)
g21828(1) = AND(g3767, g20453)
g21946(1) = AND(g5252, g18997)
g27316(1) = AND(g2407, g26710)
I24680(1) = AND(g24029, g24030, g24031, g24032)
g25921(1) = AND(g24936, g9664)
g21760(1) = AND(g3207, g20785)
g22089(1) = AND(g6311, g19210)
g28645(1) = AND(g27556, g20599)
g27342(1) = AND(g12592, g26792)
g22088(1) = AND(g6307, g19210)
g22024(1) = AND(g5897, g19147)
g27330(1) = AND(g2541, g26744)
g26099(1) = OR(g24506, g22538)
g22126(1) = AND(g6621, g19277)
g21927(1) = AND(g5164, g18997)
g23162(3) = OR(g20184, g20170, I22267)
g21755(1) = AND(g3203, g20785)
g21770(1) = AND(g3251, g20785)
g21981(1) = AND(g5543, g19074)
g22060(1) = AND(g6151, g21611)
g27087(1) = AND(g13872, g26284)
g22513(1) = NOR(g1002, g19699)
g25328(2) = AND(g5022, g23764, I24505)
g26335(1) = OR(g1526, g24609)
g21767(1) = AND(g3239, g20785)
g21794(1) = AND(g15094, g20924)
g21845(1) = AND(g3881, g21070)
g21990(1) = AND(g5591, g19074)
g21719(1) = AND(g358, g21037)
g21718(1) = AND(g370, g21037)
g21832(1) = AND(g3787, g20453)
g22055(1) = AND(g6128, g21611)
g22111(1) = AND(g6549, g19277)
g21861(1) = AND(g3949, g21070)
g24653(1) = OR(g2848, g22585)
g22070(1) = AND(g6243, g19210)
g27257(1) = OR(g25904, g24498)
g21926(1) = AND(g15147, g18997)
I24705(1) = AND(g24064, g24065, g24066, g24067)
g21701(1) = AND(g153, g20283)
g21777(1) = AND(g3380, g20391)
g22067(1) = AND(g6215, g19210)
g22094(1) = AND(g6398, g18833)
I24679(1) = AND(g19968, g24026, g24027, g24028)
g22019(1) = AND(g5857, g19147)
g22018(1) = AND(g15157, g19147)
g21997(1) = AND(g5619, g19074)
g21766(1) = AND(g3235, g20785)
g27563(1) = OR(g26104, g24704)
g27158(1) = AND(g26609, g16645)
g21871(1) = AND(g4108, g19801)
g28339(1) = AND(g9946, g27693)
g22001(1) = AND(g5731, g21562)
g22077(1) = AND(g6263, g19210)
g25848(1) = AND(g25539, g18977)
g27336(1) = AND(g2675, g26777)
g24887(2) = AND(g3712, g23239, I24054)
g21911(1) = AND(g5046, g21468)
g22102(1) = AND(g6479, g18833)
g24843(2) = AND(g3010, g23211, I24015)
g21776(1) = AND(g3376, g20391)
g21785(1) = AND(g3431, g20391)
g22066(1) = AND(g6209, g19210)
g21754(1) = AND(g3195, g20785)
I27518(1) = AND(g20720, g24104, g24105, g24106)
g27591(1) = OR(g26181, g24765)
g28315(1) = AND(g27232, g19769)
g21859(1) = AND(g3941, g21070)
g21825(1) = AND(g3736, g20453)
g21950(1) = AND(g5268, g18997)
g28257(1) = AND(g27179, g19686)
g21858(1) = AND(g3937, g21070)
g21996(1) = AND(g5615, g19074)
g21844(1) = AND(g3873, g21070)
g22076(1) = AND(g6255, g19210)
g22085(1) = AND(g6295, g19210)
g26828(1) = AND(g24919, g15756)
g22054(1) = AND(g6120, g21611)
g27580(1) = OR(g26159, g24749)
g25507(2) = AND(g6098, g23844, I24616)
I24704(1) = AND(g21193, g24061, g24062, g24063)
g21957(1) = AND(g5390, g21514)
g21739(1) = AND(g3080, g20330)
g21738(1) = AND(g3072, g20330)
g21699(1) = AND(g142, g20283)
g28706(1) = AND(g27584, g20681)
g27515(1) = OR(g26051, g13431)
g28689(1) = AND(g27575, g20651)
g28118(1) = OR(g27821, g26815)
g22131(1) = AND(g6641, g19277)
I27538(1) = AND(g21209, g24132, g24133, g24134)
g22357(1) = NOR(g1024, g19699)
g24817(1) = AND(g22929, g7235)
g26343(1) = OR(g1514, g24609)
g27294(1) = AND(g9975, g26656)
g21715(1) = AND(g160, g20283)
g22039(1) = AND(g5949, g19147)
g22038(1) = AND(g5945, g19147)
g27290(1) = OR(g25926, g25928)
g21784(1) = AND(g3423, g20391)
g21956(1) = AND(g5360, g21514)
g21889(1) = AND(g4169, g19801)
g21980(1) = AND(g5567, g19074)
g27552(1) = OR(g26092, g24676)
g21888(1) = AND(g4165, g19801)
g21824(1) = AND(g3706, g20453)
g26633(1) = AND(g24964, g20616)
g21931(1) = AND(g5188, g18997)
g22015(1) = AND(g5719, g21562)
g28269(1) = AND(g27205, g19712)
g27240(1) = OR(g25883, g24467)
g27561(1) = OR(g26100, g24702)
g22084(1) = AND(g6291, g19210)
g22110(1) = AND(g15167, g19277)
g21860(1) = AND(g3945, g21070)
g27579(1) = OR(g26157, g24748)
g21700(1) = AND(g150, g20283)
g21987(1) = AND(g5579, g19074)
g28210(1) = AND(g9229, g27554)
g21943(1) = AND(g5240, g18997)
g24558(1) = AND(g22516, g19566)
g27616(1) = AND(g26349, g20449)
g27313(1) = AND(g1982, g26701)
g21969(1) = AND(g5373, g21514)
g27276(1) = AND(g9750, g26607)
g27285(1) = AND(g9912, g26632)
g21968(1) = AND(g5459, g21514)
g27305(1) = AND(g10041, g26683)
g21855(1) = AND(g3925, g21070)
g21870(1) = AND(g4093, g19801)
g28601(1) = AND(g27506, g20514)
g27571(1) = OR(g26127, g24723)
g26329(1) = OR(g8526, g24609)
g27560(1) = AND(g26299, g20191)
g22117(1) = AND(g6597, g19277)
g22000(1) = AND(g5727, g21562)
g21867(1) = AND(g4082, g19801)
g23771(3) = OR(g21432, g21416, I22912)
g21714(1) = AND(g278, g20283)
g21707(1) = AND(g191, g20283)
g21819(1) = AND(g3614, g20924)
g21910(1) = AND(g5016, g21468)
g28666(1) = AND(g27567, g20625)
g22123(1) = AND(g6609, g19277)
g21818(1) = AND(g3610, g20924)
g21979(1) = AND(g5559, g19074)
g21978(1) = AND(g5551, g19074)
g21986(1) = AND(g5575, g19074)
g21741(1) = AND(g15086, g20330)
g21801(1) = AND(g3554, g20924)
g27974(1) = OR(g26544, g25063)
g21735(1) = AND(g3057, g20330)
g21877(1) = AND(g6888, g19801)
g22014(1) = AND(g5805, g21562)
g22007(1) = AND(g5770, g21562)
I27523(1) = AND(g20857, g24111, g24112, g24113)
g27570(1) = OR(g26126, g24722)
g22116(1) = AND(g6589, g19277)
g24984(1) = AND(g22929, g12818)
g21866(1) = AND(g4072, g19801)
g21917(1) = AND(g5092, g21468)
g22041(1) = AND(g5957, g19147)
g21706(1) = AND(g222, g20283)
g21923(1) = AND(g5029, g21468)
g22035(1) = AND(g5933, g19147)
g28587(1) = AND(g27487, g20498)
g28117(1) = AND(g8075, g27245)
g28569(1) = AND(g27453, g20433)
g22130(1) = AND(g6637, g19277)
g27284(1) = AND(g9908, g26631)
g21876(1) = AND(g4119, g19801)
g21885(1) = AND(g4122, g19801)
g27304(1) = AND(g2273, g26682)
g21854(1) = AND(g3921, g21070)
g21763(1) = AND(g3223, g20785)
g22006(1) = AND(g5767, g21562)
g27551(1) = OR(g26091, g24675)
g21916(1) = AND(g5084, g21468)
g27333(1) = AND(g10180, g26765)
g25952(1) = NOR(g1542, g24609)
g21721(1) = AND(g385, g21037)
g28586(1) = AND(g27484, g20497)
g21773(1) = AND(g3263, g20785)
g21942(1) = AND(g5236, g18997)
g22063(1) = AND(g6109, g21611)
g27312(1) = AND(g12019, g26700)
g19854(1) = NAND(I20222, I20223)
I24699(1) = AND(g21127, g24054, g24055, g24056)
I24700(1) = AND(g24057, g24058, g24059, g24060)
g23184(3) = OR(g20198, g20185, I22280)
g21734(1) = AND(g3040, g20330)
g21839(1) = AND(g3763, g20453)
g21930(1) = AND(g5180, g18997)
g21993(1) = AND(g5603, g19074)
g21838(1) = AND(g3747, g20453)
g21965(1) = AND(g15149, g21514)
I26531(1) = AND(g24099, g24100, g24101, g24102)
g25103(1) = AND(g4927, g22908)
g27184(1) = AND(g26628, g13756)
g22021(1) = AND(g5869, g19147)
g22073(1) = AND(g6235, g19210)
g27692(1) = AND(g26392, g20697)
g28193(1) = AND(g8851, g27629)
g25931(1) = AND(g24574, g19477)
g22122(1) = AND(g6601, g19277)
g22034(1) = AND(g5929, g19147)
g21815(1) = AND(g3598, g20924)
g27329(1) = AND(g12052, g26743)
g21975(1) = AND(g5523, g19074)
g27328(1) = AND(g12482, g26736)
g21937(1) = AND(g5208, g18997)
g21791(1) = AND(g3368, g20391)
g21884(1) = AND(g4104, g19801)
g27235(1) = AND(g25910, g19579)
g22109(1) = AND(g6455, g18833)
g22108(1) = AND(g6439, g18833)
g25870(1) = AND(g24840, g16182)
g25411(2) = AND(g5062, g23764, I24546)
g26094(1) = AND(g24936, g9664)
g21922(1) = AND(g5112, g21468)
g22091(1) = AND(g6415, g18833)
g21740(1) = AND(g3085, g20330)
g21953(1) = AND(g5377, g21514)
g25581(1) = AND(g19338, g24150)
g21800(1) = AND(g3546, g20924)
g21936(1) = AND(g5200, g18997)
g28346(1) = AND(g27243, g19800)
g21762(1) = AND(g3219, g20785)
g21964(1) = AND(g5441, g21514)
g23721(3) = OR(g21401, g21385, I22852)
g25067(1) = AND(g4722, g22885)
g21909(1) = AND(g5041, g21468)
g22040(1) = AND(g5953, g19147)
g27332(1) = AND(g12538, g26758)
g21908(1) = AND(g5037, g21468)
g25954(1) = NOR(g7750, g24591)
g21747(1) = AND(g3061, g20330)
g21814(1) = AND(g3594, g20924)
g21751(1) = AND(g3167, g20785)
g21807(1) = AND(g3566, g20924)
g21772(1) = AND(g3259, g20785)
g21974(1) = AND(g5517, g19074)
g22062(1) = AND(g6093, g21611)
g28108(1) = AND(g7975, g27237)
g21841(1) = AND(g3857, g21070)
g21992(1) = AND(g5599, g19074)
g25102(1) = AND(g4727, g22885)
g21835(1) = AND(g3802, g20453)
g22047(1) = AND(g6077, g21611)
g22051(1) = AND(g6105, g21611)
g22072(1) = AND(g6259, g19210)
g28192(1) = AND(g8891, g27415)
g21720(1) = AND(g376, g21037)
g28663(1) = AND(g27566, g20624)
g21746(1) = AND(g3045, g20330)
g21983(1) = AND(g5555, g19074)
g21806(1) = AND(g3558, g20924)
g27325(1) = AND(g12478, g26724)
g25085(1) = AND(g4912, g22908)
g22020(1) = AND(g5863, g19147)
g27291(1) = AND(g11969, g26653)
g22046(1) = AND(g6073, g21611)
g22113(1) = AND(g6561, g19277)
g21863(1) = AND(g3957, g21070)
g26327(1) = OR(g8462, g24591)
g22105(1) = AND(g6494, g18833)
g26342(1) = OR(g8407, g24591)
g21703(1) = AND(g146, g20283)
g21781(1) = AND(g3408, g20391)
g21952(1) = AND(g5366, g21514)
g28311(1) = AND(g9792, g27679)
g21821(1) = AND(g3723, g20453)
g21790(1) = AND(g3454, g20391)
g21873(1) = AND(g6946, g19801)
g22027(1) = AND(g5889, g19147)
g21834(1) = AND(g3752, g20453)
g22003(1) = AND(g5736, g21562)
g26084(1) = AND(g24926, g9602)
g25143(1) = AND(g4922, g22908)
g22081(1) = AND(g6279, g19210)
g27633(1) = AND(g13076, g25766)
g21913(1) = AND(g5069, g21468)
g25479(1) = AND(g22646, g9917)
g22090(1) = AND(g6404, g18833)
g27247(1) = AND(g2759, g26745)
g21797(1) = AND(g3518, g20924)
g25580(1) = AND(g19268, g24149)
g22523(1) = NOR(g1345, g19720)
g28113(1) = AND(g8016, g27242)
g27099(1) = AND(g14094, g26352)
g27324(1) = AND(g10150, g26720)
g25084(1) = AND(g4737, g22885)
g22026(1) = AND(g5913, g19147)
g25417(2) = AND(g5712, g23816, I24552)
g21711(1) = AND(g291, g20283)
g22097(1) = AND(g6451, g18833)
g22104(1) = AND(g6444, g18833)
g21750(1) = AND(g3161, g20785)
g28248(1) = AND(g27150, g19676)
g27589(1) = OR(g26177, g24763)
g21982(1) = AND(g5547, g19074)
g21796(1) = AND(g3512, g20924)
g24782(3) = OR(g23857, g23872)
g22133(1) = AND(g6649, g19277)
I24685(1) = AND(g24036, g24037, g24038, g24039)
g21840(1) = AND(g15099, g21070)
g22011(1) = AND(g15154, g21562)
g25123(1) = AND(g4732, g22885)
g24578(1) = OR(g2882, g23825)
g22112(1) = AND(g6555, g19277)
g21862(1) = AND(g3953, g21070)
g22050(1) = AND(g6088, g21611)
g21949(1) = AND(g5264, g18997)
g21948(1) = AND(g5260, g18997)
g22096(1) = AND(g6434, g18833)
g21702(1) = AND(g157, g20283)
g21757(1) = AND(g3187, g20785)
g25579(1) = AND(g19422, g24147)
g25578(1) = AND(g19402, g24146)
g26334(1) = OR(g1171, g24591)
g22539(1) = NOR(g1030, g19699)
g24890(1) = NAND(g13852, g22929)
g21847(1) = AND(g3905, g21070)
g27281(1) = AND(g9830, g26615)
g21933(1) = AND(g5212, g18997)
g27301(1) = AND(g11992, g26679)
g25947(1) = NOR(g1199, g24591)
g21851(1) = AND(g3901, g21070)
g21872(1) = AND(g4098, g19801)
g27699(1) = AND(g26396, g20766)
g22129(1) = AND(g6633, g19277)
g22002(1) = AND(g5706, g21562)
g22057(1) = AND(g15159, g21611)
g22128(1) = AND(g6629, g19277)
g25142(1) = AND(g4717, g22885)
g21912(1) = AND(g5052, g21468)
g26821(1) = AND(g24821, g13103)
g21756(1) = AND(g3211, g20785)
g21780(1) = AND(g3391, g20391)
g28369(1) = OR(g27160, g25938)
g21820(1) = AND(g3712, g20453)
g28627(1) = AND(g27543, g20574)
g21846(1) = AND(g3897, g21070)
g21731(1) = AND(g3029, g20330)
g21929(1) = AND(g5176, g18997)
g22056(1) = AND(g6133, g21611)
g21928(1) = AND(g5170, g18997)
g22080(1) = AND(g6275, g19210)
g24858(2) = AND(g3361, g23223, I24030)
g25873(1) = AND(g24854, g16197)
g21787(1) = AND(g15091, g20391)
g22031(1) = AND(g5917, g19147)
g21743(1) = AND(g3100, g20330)
g21827(1) = AND(g3759, g20453)
g21769(1) = AND(g3247, g20785)
g25453(2) = AND(g5406, g23789, I24576)
g21768(1) = AND(g3243, g20785)
g21803(1) = AND(g3538, g20924)
g28299(1) = AND(g9716, g27670)
g22132(1) = AND(g6645, g19277)
g21881(1) = AND(g4064, g19801)
g22491(1) = NOR(g1361, g19720)
g25905(1) = AND(g24879, g16311)
g22087(1) = AND(g6303, g19210)
g21890(1) = AND(g4125, g19801)
g25958(1) = NOR(g7779, g24609)
g27581(1) = OR(g26161, g24750)
g22043(1) = AND(g5965, g19147)
g21710(1) = AND(g287, g20283)
g21779(1) = AND(g3385, g20391)
g26750(1) = AND(g24514, g24474)
g22069(1) = AND(g6227, g19210)
g25408(1) = AND(g22682, g9772)
g21778(1) = AND(g3355, g20391)
g22068(1) = AND(g6219, g19210)
g21786(1) = AND(g3436, g20391)
g21945(1) = AND(g5248, g18997)
g21826(1) = AND(g3742, g20453)
g21999(1) = AND(g5723, g21562)
g27315(1) = AND(g12022, g26709)
g21998(1) = AND(g5712, g21562)
g21932(1) = AND(g5204, g18997)
g22010(1) = AND(g5787, g21562)
g21961(1) = AND(g5424, g21514)
g22079(1) = AND(g6271, g19210)
g22078(1) = AND(g6267, g19210)
g21717(1) = AND(g15051, g21037)
g22086(1) = AND(g6299, g19210)
g28330(1) = AND(g27238, g19786)
g22125(1) = AND(g6617, g19277)
g21811(1) = AND(g3582, g20924)
g28258(1) = AND(g27182, g19687)
g21971(1) = AND(g5417, g21514)
g27256(1) = AND(g25937, g19698)
g22017(1) = AND(g5763, g21562)
g27280(1) = AND(g9825, g26614)
g27300(1) = AND(g12370, g26672)
g21850(1) = AND(g3893, g21070)
g28602(1) = AND(g27509, g20515)
g27562(1) = OR(g26102, g24703)
g22023(1) = AND(g5881, g19147)
g21716(1) = AND(g301, g20283)
g21959(1) = AND(g5413, g21514)
g21925(1) = AND(g5073, g21468)
g28919(1) = AND(g27663, g21295)
g21958(1) = AND(g5396, g21514)
g21742(1) = AND(g3050, g20330)
g21944(1) = AND(g5244, g18997)
g27314(1) = AND(g12436, g26702)
g21802(1) = AND(g3562, g20924)
g21857(1) = AND(g3933, g21070)
g21730(1) = AND(g3025, g20330)
g21793(1) = AND(g3412, g20391)
g28159(1) = AND(g8553, g27317)
g22016(1) = AND(g5747, g21562)
g27394(1) = OR(g25957, g24573)
g21765(1) = AND(g3231, g20785)
g27341(1) = AND(g10203, g26788)
g27335(1) = AND(g12087, g26776)
g22042(1) = AND(g5961, g19147)
g27667(1) = AND(g26361, g20601)
g22124(1) = AND(g6613, g19277)
g22030(1) = AND(g5909, g19147)
g19782(1) = NAND(I20188, I20189)
g22093(1) = AND(g6423, g18833)
g21775(1) = AND(g3372, g20391)
g22065(1) = AND(g6203, g19210)
g21737(1) = AND(g3068, g20330)
g27286(1) = AND(g6856, g26634)
g21856(1) = AND(g3929, g21070)
g21995(1) = AND(g5611, g19074)
g21880(1) = AND(g4135, g19801)
g27677(1) = AND(g13021, g25888)
g26779(1) = AND(g24497, g23620)
g21831(1) = AND(g3782, g20453)
I25736(1) = OR(g12, g22150, g20277)
g22535(1) = NOR(g19699, g1030)
g24018(1) = NOR(I23162, I23163)
g24965(1) = OR(g22667, g23825)
g24468(2) = OR(g10925, g22400)
g22540(1) = NOR(g19720, g1373)
g24363(1) = OR(g7831, g22138)
g24478(2) = OR(g11003, g22450)
g24433(2) = OR(g10878, g22400)
g24460(2) = OR(g10967, g22450)
g24661(1) = NAND(g23210, g23195, g22984)
g24620(1) = NAND(g22902, g22874)
g22488(1) = NOR(g19699, g1002)
g22537(1) = NOR(g19720, g1367)
g24566(1) = NAND(g22755, g22713)
g24678(1) = NAND(g22994, g23010)
g22522(1) = NOR(g19699, g1024)
g25010(1) = OR(g23267, g2932)
g24880(1) = NAND(g23281, g23266, g22839)
g24447(2) = OR(g10948, g22450)
g24544(1) = NAND(g22666, g22661, g22651)
g24547(1) = NAND(g22638, g22643, g22754)
g24652(1) = NAND(g22712, g22940, g22757)
g24457(2) = OR(g10902, g22400)
g24471(2) = OR(g10999, g22450)
g24444(2) = OR(g10890, g22400)
g22514(1) = NOR(g19699, g1018)
g22517(1) = NOR(g19720, g1345)
g24584(1) = NAND(g22852, g22836, g22715)
g22524(1) = NOR(g19720, g1361)
I22761(1) = NAND(g11939, I22760)
g24362(1) = NAND(g21370, g22136)
I22973(1) = NAND(g9657, I22972)
I22974(1) = NAND(g19638, I22972)
I22800(1) = NAND(g11960, I22799)
I22801(1) = NAND(g21434, I22799)
I22946(1) = NAND(g19620, I22944)
I22755(1) = NAND(g21434, I22753)
I22794(1) = NAND(g21434, I22792)
I22845(1) = NAND(g12113, I22844)
I22762(1) = NAND(g21434, I22760)
I22719(1) = NAND(g21434, I22717)
I22718(1) = NAND(g11916, I22717)
I22754(1) = NAND(g11937, I22753)
I22872(1) = NAND(g12150, I22871)
I22873(1) = NAND(g21228, I22871)
I22966(1) = NAND(g12288, I22965)
I22967(1) = NAND(g21228, I22965)
I22824(1) = NAND(g21434, I22822)
I22931(1) = NAND(g21228, I22929)
I22893(1) = NAND(g12189, I22892)
I22894(1) = NAND(g21228, I22892)
I22866(1) = NAND(g21228, I22864)
I22921(2) = NAND(g14677, g21284)
I22930(1) = NAND(g12223, I22929)
I22937(1) = NAND(g12226, I22936)
I22685(1) = NAND(g21434, I22683)
I22846(1) = NAND(g21228, I22844)
I21978(1) = NAND(g19620, I21976)
g23975(3) = NAND(I23119, I23120)
I22684(1) = NAND(g11893, I22683)
I21993(1) = NAND(g7670, I21992)
I22711(1) = NAND(g11915, I22710)
I22793(1) = NAND(g11956, I22792)
I22945(1) = NAND(g9492, I22944)
I22823(1) = NAND(g11978, I22822)
I21977(1) = NAND(g7680, I21976)
I22900(1) = NAND(g12193, I22899)
I22901(1) = NAND(g21228, I22899)
I22865(1) = NAND(g12146, I22864)
I22938(1) = NAND(g21228, I22936)
I22712(1) = NAND(g21434, I22710)
g27377(1) = NAND(g10685, g25930)
I21994(1) = NAND(g19638, I21992)
g23002(1) = NOT(I22177)
g23612(1) = NOT(I22745)
g23652(1) = NOT(I22785)
g23759(1) = NOT(I22886)
g25582(1) = OR(g21662, g24152)
g25583(1) = OR(g21666, g24153)
g25584(1) = OR(g21670, g24154)
g25585(1) = OR(g21674, g24155)
g25586(1) = OR(g21678, g24156)
g25587(1) = OR(g21682, g24157)
g25588(1) = OR(g21686, g24158)
g25589(1) = OR(g21690, g24159)
g25590(1) = OR(g21694, g24160)
g29301(1) = OR(g28686, g18797)
g28051(1) = OR(g27699, g18166)
g29282(1) = OR(g28617, g18745)
g26920(1) = OR(g25865, g18283)
g29296(1) = OR(g28586, g18781)
g28047(1) = OR(g27676, g18160)
g29273(1) = OR(g28269, g18639)
g29265(1) = OR(g28318, g18620)
g29295(1) = OR(g28663, g18780)
g29306(1) = OR(g28689, g18813)
g29272(1) = OR(g28346, g18638)
g29283(1) = OR(g28627, g18746)
g29224(1) = OR(g28919, g18156)
g28052(1) = OR(g27710, g18167)
g29294(1) = OR(g28645, g18779)
g28050(1) = OR(g27692, g18165)
g29293(1) = OR(g28570, g18777)
g29264(1) = OR(g28248, g18618)
g29271(1) = OR(g28333, g18637)
g29261(1) = OR(g28247, g18605)
g28055(1) = OR(g27560, g18190)
g29307(1) = OR(g28706, g18814)
g29270(1) = OR(g28258, g18635)
g26926(1) = OR(g26633, g18531)
g29266(1) = OR(g28330, g18621)
g28060(1) = OR(g27616, g18532)
g29300(1) = OR(g28666, g18796)
g28058(1) = OR(g27235, g18268)
g29267(1) = OR(g28257, g18622)
g25623(1) = OR(g24552, g18219)
g29305(1) = OR(g28602, g18811)
g29302(1) = OR(g28601, g18798)
g29290(1) = OR(g28569, g18764)
g29287(1) = OR(g28555, g18760)
g28046(1) = OR(g27667, g18157)
g29289(1) = OR(g28642, g18763)
g29281(1) = OR(g28541, g18743)
g28049(1) = OR(g27684, g18164)
g26913(1) = OR(g25848, g18225)
g28044(1) = OR(g27256, g18130)
g26925(1) = OR(g25939, g18301)
g29299(1) = OR(g28587, g18794)
g29284(1) = OR(g28554, g18747)
g29288(1) = OR(g28630, g18762)
g26918(1) = OR(g25931, g18243)
g28056(1) = OR(g27230, g18210)
g29308(1) = OR(g28612, g18815)
g29260(1) = OR(g28315, g18604)
g25632(1) = OR(g24558, g18277)
g29259(1) = OR(g28304, g18603)
g28054(1) = OR(g27723, g18170)
g29258(1) = OR(g28238, g18601)
I24041(1) = NOT(g22182)
I24191(1) = NOT(g22360)
g23823(1) = NOT(I22989)
g22228(69) = NOT(I21810)
g23650(1) = NOT(g20653)
g22594(27) = NOT(I21934)
g26673(5) = OR(g24433, g10674)
g23529(1) = NOT(g20558)
g24518(3) = OR(g22517, g7601)
g28431(3) = NOT(I26925)
g25356(1) = NOT(g22763)
g22722(28) = NOT(I22031)
g23776(1) = NOT(g21177)
g25182(1) = NOT(g22763)
I23384(1) = NOT(g23362)
g23870(1) = NOT(g21293)
I24781(1) = NOT(g24264)
g25212(1) = NOT(g22763)
g27662(1) = NOT(I26296)
I23351(1) = NOT(g23263)
I23348(1) = NOT(g23384)
g25011(1) = NOT(g22763)
g28353(3) = NOR(g9073, g27654, g24732)
g26725(5) = OR(g24457, g10719)
I23381(1) = NOT(g23322)
I23378(1) = NOT(g23426)
I24474(1) = NOT(g22546)
g22171(1) = NOT(g18882)
g25549(1) = NOT(g22763)
g22550(34) = NOT(I21922)
g25245(1) = NOT(g22763)
g25299(1) = NOT(g22763)
g23760(1) = NOT(I22889)
I23333(1) = NOT(g22683)
g25316(1) = NOT(g22763)
g25529(1) = NOT(g22763)
g26337(1) = NOT(g24818)
I23339(1) = NOT(g23232)
I24445(1) = NOT(g22923)
g24537(2) = AND(g22626, g10851)
I23369(1) = NOT(g23347)
I24787(1) = NOT(g24266)
I24497(1) = NOT(g22592)
I23345(1) = NOT(g23320)
I23399(1) = NOT(g23450)
g25531(1) = NAND(g22763, g2868)
I23336(1) = NOT(g22721)
g23231(1) = NOT(g20050)
g25224(1) = NOT(g22763)
I25356(1) = NOT(g24374)
g25308(1) = NOT(g22763)
I24331(1) = NOT(g22976)
I24448(1) = NOT(g22923)
g24982(1) = NOT(g22763)
I23366(1) = NOT(g23321)
g25195(1) = NOT(g22763)
g23800(1) = NOT(g21246)
g24485(2) = AND(g10710, g22319)
g24541(2) = AND(g22626, g10851)
g29190(1) = NOT(g27046)
g23653(1) = NOT(I22788)
I23688(1) = NOT(g23244)
I24228(1) = NOT(g22409)
I23393(1) = NOT(g23414)
g23745(1) = NOT(g20900)
g28325(1) = NOT(g27463)
g27093(1) = NOR(g26712, g26749)
g28504(3) = NAND(g758, g27528, g11679)
g24756(1) = NOT(g22763)
g25194(1) = NOT(g22763)
g29196(1) = NOT(g27059)
I22819(1) = NOT(g19862)
I22816(1) = NOT(g19862)
g29933(3) = NOR(g8808, g28500, g12259)
g28444(3) = NOR(g8575, g27463, g24825)
g26818(1) = NOT(I25530)
I23360(1) = NOT(g23360)
g26793(5) = OR(g24478, g7520)
I23390(1) = NOT(g23395)
g23613(1) = NOT(I22748)
g25438(1) = NOT(g22763)
g25348(1) = NOT(g22763)
g28370(1) = NOT(g27528)
I24078(1) = NOT(g22360)
g24715(1) = OR(g22189, g22207)
I24022(1) = NOT(g22182)
g26759(5) = OR(g24468, g7511)
g30184(1) = NOT(g28144)
I23354(1) = NOT(g23277)
g25184(1) = NOT(g22763)
I23671(1) = NOT(g23202)
g27102(1) = NOR(g26750, g26779)
g23651(1) = NOT(g20655)
g23440(2) = NOT(I22557)
g25882(1) = NOT(g25026)
g24995(1) = NOT(g22763)
g24491(2) = AND(g10727, g22332)
g25399(1) = NOT(g22763)
I24455(1) = NOT(g22541)
g25263(1) = NOT(g22763)
I23327(1) = NOT(g22647)
g26703(5) = OR(g24447, g10705)
I23357(1) = NOT(g23359)
g25541(1) = NOT(g22763)
g25535(1) = NOT(g22763)
I24008(1) = NOT(g22182)
g23715(1) = NOT(g20764)
I23694(1) = NOT(g23252)
g24966(1) = NOT(g22763)
g23824(1) = NOT(g21271)
I25190(1) = NOT(g25423)
g26737(5) = OR(g24460, g10720)
I24215(1) = NOT(g22360)
g25262(1) = NOT(g22763)
g25899(1) = NOT(g24997)
I23363(1) = NOT(g23385)
I24060(1) = NOT(g22202)
g25388(1) = NOT(g22763)
g25534(1) = NOT(g22763)
g26770(5) = OR(g24471, g10732)
g28479(1) = NOT(g27654)
g25227(1) = NOT(g22763)
I23680(1) = NOT(g23219)
g25562(1) = NOT(g22763)
g27585(1) = NOT(g25994)
I23684(1) = NOT(g23230)
I23375(1) = NOT(g23403)
g27576(1) = NOT(g26081)
I23342(1) = NOT(g23299)
g25226(1) = NOT(g22763)
g23746(1) = NOT(g20902)
I23372(1) = NOT(g23361)
g25211(1) = NOT(g22763)
I24434(1) = NOT(g22763)
g28137(1) = NOT(I26638)
g28174(3) = NAND(g1270, g27059)
I23396(1) = NOT(g23427)
g25196(1) = NOT(g22763)
g25537(1) = NAND(g22763, g2873)
g25550(1) = NOT(g22763)
g25307(1) = NOT(g22763)
g23003(1) = NOT(I22180)
g25243(1) = NOT(g22763)
g24744(2) = NOT(g22202)
I26989(1) = NOT(g27277)
g25557(1) = NOT(g22763)
g28314(1) = AND(g27552, g14205)
I22576(1) = NOT(g21282)
g25169(1) = NOT(g22763)
I24334(1) = NOT(g22976)
g25556(1) = NOT(g22763)
I24089(1) = NOT(g22409)
I23998(1) = NOT(g22182)
g24641(1) = OR(g22151, g22159)
I24784(1) = NOT(g24265)
I23387(1) = NOT(g23394)
g24770(1) = NOT(g22763)
g24981(1) = NOT(g22763)
g24718(2) = NOT(g22182)
g25340(1) = NOT(g22763)
g25193(1) = NOT(g22763)
I23330(1) = NOT(g22658)
g24510(3) = OR(g22488, g7567)
g24996(1) = NOT(g22763)
g25209(1) = NOT(g22763)
g26694(5) = OR(g24444, g10704)
g25208(1) = NOT(g22763)
g25542(1) = NOT(g22763)
g25274(1) = NOT(g22763)
g25283(1) = NOT(g22763)
g24872(2) = AND(g23088, g9104)
I24038(1) = NOT(g22202)
g25183(1) = NOT(g22763)
g28167(3) = NAND(g925, g27046)
g28598(1) = NOT(g27717)
g29745(1) = NOT(g28500)
g25282(1) = NOT(g22763)
g25768(1) = AND(g2912, g24560)
g28558(1) = AND(g7301, g27046)
g28679(1) = AND(g27572, g20638)
g27964(1) = AND(g25956, g22492)
g25331(2) = AND(g5366, g22194, I24508)
g28160(1) = AND(g26309, g27463)
g28605(1) = OR(g27341, g26302)
g28455(1) = AND(g27289, g20103)
g23616(1) = NAND(I22754, I22755)
g25149(1) = AND(g14030, g23546)
g25148(1) = AND(g16867, g23545)
g28591(1) = OR(g27332, g26286)
g25104(1) = AND(g16800, g23504)
g23748(1) = NAND(I22872, I22873)
g26785(2) = OR(g10776, g24468)
g25850(1) = AND(g3502, g24636)
g24884(2) = AND(g3401, g23555, I24051)
g28566(1) = OR(g27316, g26254)
g25062(1) = NAND(g21403, g23363)
g25049(1) = NAND(g21344, g23462)
g24666(1) = AND(g11753, g22975)
g28546(1) = OR(g27302, g26231)
g27532(1) = OR(g16176, g26084)
g27231(1) = OR(g25873, g15699)
g26789(2) = OR(g10776, g24471)
g28285(1) = AND(g9657, g27717)
g25112(1) = AND(g10428, g23510)
g27035(1) = AND(g26348, g1500)
g24654(1) = AND(g11735, g22922)
g24989(1) = NAND(g21345, g23363)
g24973(1) = NAND(g21272, g23462)
g27362(1) = AND(g26080, g20036)
g28712(1) = AND(g27590, g20708)
g25129(1) = AND(g17682, g23527)
g25128(1) = AND(g17418, g23525)
g26755(2) = OR(g10776, g24457)
g27026(1) = OR(g26828, g17726)
g25775(1) = AND(g2922, g24568)
g24772(1) = AND(g16287, g23061)
g24638(1) = AND(g22763, g19690)
g25831(1) = AND(g3151, g24623)
g24835(1) = AND(g8720, g23233)
g28603(1) = OR(g27340, g26300)
g25056(1) = AND(g12779, g23456)
g27034(1) = AND(g26328, g8609)
g28653(1) = AND(g7544, g27014)
g29078(1) = OR(g27633, g26572)
g25031(1) = AND(g20675, g23432)
g28614(1) = OR(g27351, g26311)
g27250(1) = OR(g25901, g15738)
g24684(1) = AND(g11769, g22989)
g25132(1) = AND(g10497, g23528)
g25087(1) = AND(g17307, g23489)
g24727(1) = AND(g13300, g23016)
g25043(1) = AND(g20733, g23447)
g26079(1) = AND(g6199, g25060)
g28674(1) = AND(g27569, g20629)
g25068(1) = AND(g17574, g23477)
g28526(1) = OR(g27285, g26178)
g28692(1) = AND(g27578, g20661)
g28536(1) = OR(g27293, g26205)
g28581(1) = OR(g27329, g26276)
g28613(1) = OR(g27350, g26310)
g25079(1) = AND(g21011, g23483)
g25086(1) = AND(g13941, g23488)
g24726(1) = AND(g15965, g23015)
g26733(2) = OR(g10776, g24447)
g25125(1) = AND(g20187, g23520)
g26805(2) = OR(g10776, g24478)
g24635(1) = AND(g19874, g22883)
g26842(1) = AND(g2894, g24522)
g28725(1) = AND(g27596, g20779)
g25571(1) = AND(I24694, I24695)
g28107(1) = AND(g27970, g18874)
g23747(1) = NAND(I22865, I22866)
g22920(1) = AND(g19764, g19719)
g26294(1) = AND(g4245, g25230)
g28580(1) = OR(g27328, g26275)
g24663(1) = AND(g16621, g22974)
g24949(1) = AND(g23796, g20751)
g24536(1) = AND(g19516, g22635)
g24904(1) = AND(g11761, g23279)
g25093(1) = AND(g12831, g23493)
g24564(1) = AND(g23198, g21163)
g28525(1) = OR(g27284, g26176)
g26853(1) = AND(g94, g24533)
g25201(1) = AND(g12346, g23665)
g24912(1) = AND(g23687, g20682)
g26864(1) = AND(g2907, g24548)
g25782(1) = AND(g2936, g24571)
g23655(1) = NAND(I22793, I22794)
g22861(1) = AND(g19792, g19670)
g26344(1) = OR(g2927, g25010)
g27932(1) = AND(g25944, g19369)
g28574(1) = OR(g27324, g26270)
g24846(2) = AND(g3361, g23555, I24018)
g28551(1) = OR(g27305, g26234)
g24929(1) = AND(g23751, g20875)
g28517(1) = OR(g27280, g26154)
g24968(2) = OR(g22360, g22409, g23389)
g27097(1) = AND(g25867, g22526)
g25894(1) = OR(g24817, g23229)
g24769(1) = AND(g19619, g23058)
g25166(1) = AND(g17506, g23571)
g27274(1) = OR(g15779, g25915)
g28573(1) = AND(g7349, g27059)
g25485(2) = AND(g6098, g22220, I24600)
g25570(1) = AND(I24689, I24690)
g27959(1) = AND(g25948, g19374)
g27050(1) = AND(g25789, g22338)
g27958(1) = AND(g25950, g22449)
g25907(1) = AND(g24799, g22519)
g25567(1) = AND(I24674, I24675)
g25238(1) = AND(g12466, g23732)
g24647(1) = AND(g19903, g22907)
g26304(1) = AND(g2697, g25246)
g24998(1) = AND(g17412, g23408)
g24672(1) = AND(g19534, g22981)
g28533(1) = OR(g27291, g26203)
g28451(1) = AND(g27283, g20090)
g24975(1) = NAND(g21388, g23363)
g24958(1) = NAND(g21330, g23462)
g28596(1) = OR(g27336, g26291)
g27323(1) = AND(g26268, g23086)
g28595(1) = OR(g27335, g26290)
g24946(2) = OR(g22360, g22409, g8130)
g26312(1) = AND(g2704, g25264)
g29325(1) = OR(g28813, g27820)
g24716(1) = AND(g15935, g23004)
g27224(1) = OR(g25870, g15678)
g24627(1) = AND(g22763, g19679)
g23780(1) = NAND(I22930, I22931)
g27393(1) = AND(g26099, g20066)
g27258(1) = OR(g25905, g15749)
g24681(1) = AND(g16653, g22988)
g24549(1) = AND(g23162, g20887)
g25207(1) = AND(g22513, g10621)
g27043(1) = AND(g26335, g8632)
g28426(1) = AND(g27257, g20006)
g26849(1) = AND(g2994, g24527)
g25414(2) = AND(g5406, g22194, I24549)
g26848(1) = AND(g2950, g24526)
g28560(1) = OR(g27311, g26249)
g27086(1) = AND(g25836, g22495)
g26833(1) = AND(g2852, g24509)
g28658(1) = AND(g27563, g20611)
g25107(1) = AND(g17643, g23508)
g26048(1) = AND(g5853, g25044)
g28592(1) = OR(g27333, g26288)
g28279(1) = OR(g27087, g25909)
g28714(1) = AND(g27591, g20711)
g24709(1) = AND(g16690, g23000)
g24708(1) = AND(g16474, g22998)
g29475(1) = AND(g14033, g28500)
g25106(1) = AND(g17391, g23506)
g24602(1) = AND(g16507, g22854)
g25033(1) = AND(g17500, g23433)
g25371(2) = AND(g5062, g22173, I24524)
g26829(1) = AND(g2844, g24505)
g26766(2) = OR(g10776, g24460)
g28695(1) = AND(g27580, g20666)
g23576(1) = NAND(I22718, I22719)
g25163(1) = AND(g20217, g23566)
g28577(1) = OR(g27326, g26272)
g25012(1) = AND(g20644, g23419)
g28597(1) = AND(g27515, g20508)
g30173(1) = AND(g28118, g13082)
g23761(1) = NAND(I22893, I22894)
g28368(1) = OR(g27158, g27184)
g25960(1) = OR(g24566, g24678)
g27030(1) = AND(g26343, g7947)
g24656(1) = AND(g11736, g22926)
g25173(1) = AND(g12234, g23589)
g24680(1) = AND(g16422, g22986)
g28456(1) = AND(g27290, g20104)
g28341(1) = AND(g27240, g19790)
g29643(1) = OR(g28192, g27145)
g25021(1) = NAND(g21417, g23363)
g25003(1) = NAND(g21353, g23462)
g28655(1) = AND(g27561, g20603)
g28694(1) = AND(g27579, g20664)
g23656(1) = NAND(I22800, I22801)
g26690(2) = OR(g10776, g24433)
g24668(1) = AND(g11754, g22979)
g28549(1) = OR(g27304, g26233)
g27119(1) = AND(g25877, g22542)
g28548(1) = OR(g27303, g26232)
g25038(1) = NAND(g21331, g23363)
g25020(1) = NAND(g21377, g23462)
g25573(1) = AND(I24704, I24705)
g24865(1) = AND(g11323, g23253)
g25045(1) = AND(g17525, g23448)
g28677(1) = AND(g27571, g20635)
g27036(1) = AND(g26329, g11038)
g24679(1) = AND(g13289, g22985)
g23575(1) = NAND(I22711, I22712)
g25462(2) = AND(g6404, g22300, I24585)
g24939(1) = AND(g23771, g21012)
g25061(1) = AND(g17586, g23461)
g26858(1) = AND(g2970, g24540)
g28110(1) = AND(g27974, g18886)
g28607(1) = OR(g27342, g26303)
g28625(1) = OR(g27363, g26324)
g26721(2) = OR(g10776, g24444)
g27019(1) = OR(g26822, g14610)
g25071(1) = AND(g12804, g23478)
g28676(1) = AND(g27570, g20632)
g25147(1) = AND(g20202, g23542)
g25151(1) = AND(g17719, g23549)
g26301(1) = AND(g2145, g25244)
g24822(2) = AND(g3010, g23534, I24003)
g25420(2) = AND(g6058, g22220, I24555)
g28576(1) = OR(g27325, g26271)
g25059(1) = AND(g20870, g23460)
g27083(1) = AND(g25819, g22456)
g24864(1) = AND(g11201, g22305)
g25377(2) = AND(g5712, g22210, I24530)
g24900(2) = AND(g3752, g23582, I24067)
g28638(1) = AND(g27551, g20583)
g25290(2) = AND(g5022, g22173, I24482)
g24642(1) = AND(g8290, g22898)
g27963(1) = AND(g25952, g16047)
g27278(1) = OR(g15786, g25921)
g28545(1) = OR(g27301, g26230)
g24892(1) = AND(g11559, g23264)
g24476(1) = AND(g18879, g22330)
g22873(1) = AND(g19854, g19683)
g25572(1) = AND(I24699, I24700)
g29319(1) = OR(g28812, g14453)
g24555(1) = AND(g23184, g21024)
g24712(1) = AND(g19592, g23001)
g24914(1) = AND(g8721, g23301)
g25127(1) = AND(g13997, g23524)
g28237(1) = AND(g9492, g27597)
g26088(1) = AND(g6545, g25080)
g28538(1) = OR(g27294, g26206)
g24637(1) = AND(g16586, g22884)
g28165(1) = AND(g27018, g22455)
g28582(1) = OR(g27330, g26277)
g26855(1) = AND(g2960, g24535)
g28448(2) = NAND(g23975, g27377)
g24729(1) = AND(g22719, g23018)
g25088(1) = AND(g17601, g23491)
g24728(1) = AND(g16513, g23017)
g23719(1) = NAND(I22845, I22846)
g25126(1) = AND(g16839, g23523)
g24622(1) = AND(g19856, g22866)
g26257(1) = AND(g4253, g25197)
g28565(1) = OR(g27315, g26253)
g26019(1) = AND(g5507, g25032)
g28544(1) = OR(g27300, g26229)
g25986(1) = AND(g5160, g25013)
g24921(1) = AND(g23721, g20739)
g23781(1) = NAND(I22937, I22938)
g25150(1) = AND(g17480, g23547)
g27962(1) = AND(g25954, g19597)
g28164(1) = AND(g8651, g27528)
g26854(1) = AND(g2868, g24534)
g25866(1) = AND(g3853, g24648)
g28518(1) = OR(g27281, g26158)
g26287(1) = AND(g2138, g25225)
g26839(1) = AND(g2988, g24516)
g25456(2) = AND(g5752, g22210, I24579)
g26838(1) = AND(g2860, g24515)
g25076(1) = AND(g12805, g23479)
g25054(1) = AND(g12778, g23452)
g24725(1) = AND(g19587, g23012)
g26279(1) = AND(g4249, g25213)
g28589(1) = OR(g27331, g26285)
g27024(1) = OR(g26826, g17692)
g24849(1) = AND(g4165, g22227)
g26363(1) = OR(g2965, g24965)
g27029(1) = AND(g26327, g11031)
g27028(1) = AND(g26342, g1157)
g29114(1) = OR(g27646, g26602)
g25187(1) = AND(g12296, g23629)
g28152(1) = AND(g26297, g27279)
g24812(1) = AND(g19662, g22192)
g26186(1) = AND(g24580, g23031)
g28534(1) = OR(g27292, g26204)
g28564(1) = OR(g27314, g26252)
g25217(1) = AND(g12418, g23698)
g25223(1) = AND(g22523, g10652)
g25887(1) = NOR(g24984, g11706)
g23762(1) = NAND(I22900, I22901)
g27098(1) = AND(g25868, g22528)
g23809(1) = NAND(I22966, I22967)
g25110(1) = AND(g10427, g23509)
g24788(1) = AND(g11384, g23111)
g25179(1) = AND(g16928, g23611)
g25178(1) = AND(g20241, g23608)
g27140(1) = AND(g25885, g22593)
g23685(1) = NAND(I22823, I22824)
g23617(1) = NAND(I22761, I22762)
g28710(1) = AND(g27589, g20703)
g28204(1) = AND(g26098, g27654)
g25908(1) = AND(g24782, g22520)
g25569(1) = AND(I24684, I24685)
g25568(1) = AND(I24679, I24680)
g28182(1) = AND(g8770, g27349)
g24944(1) = NAND(g21354, g23363)
g24934(1) = NAND(g21283, g23462)
g28672(1) = AND(g7577, g27017)
g24755(1) = AND(g16022, g23030)
g24794(1) = AND(g11414, g23138)
g25510(2) = AND(g6444, g22300, I24619)
g27025(1) = AND(g26334, g7917)
g25014(1) = AND(g17474, g23420)
g28527(1) = OR(g27286, g26182)
g26130(1) = AND(g24890, g19772)
g24861(2) = AND(g3712, g23582, I24033)
g27957(1) = AND(g25947, g15995)
g27120(1) = AND(g25878, g22543)
g24974(1) = NAND(g21301, g23363)
g24957(1) = NAND(g21359, g23462)
g24777(1) = AND(g11345, g23066)
g23552(1) = NAND(I22684, I22685)
g25165(1) = AND(g14062, g23570)
g29837(1) = AND(g28369, g20144)
g28594(1) = OR(g27334, g26289)
g24754(1) = AND(g19604, g23027)
g26274(1) = AND(g2130, g25210)
g26292(1) = AND(g2689, g25228)
g28578(1) = OR(g27327, g26273)
g27542(1) = OR(g16190, g26094)
g29477(1) = AND(g14090, g28441)
g27968(1) = AND(g25958, g19614)
g28697(1) = AND(g27581, g20669)
g28562(1) = OR(g27313, g26251)
g28561(1) = OR(g27312, g26250)
g25164(1) = AND(g16883, g23569)
g28198(1) = AND(g26649, g27492)
g25091(1) = AND(g12830, g23492)
g25192(1) = AND(g20276, g23648)
g26847(1) = AND(g2873, g24525)
g25040(1) = AND(g12738, g23443)
g28657(1) = AND(g27562, g20606)
g27016(1) = OR(g26821, g14585)
g24644(1) = AND(g11714, g22903)
g24855(2) = AND(g3050, g23534, I24027)
g28513(1) = OR(g27276, g26123)
g26846(1) = AND(g37, g24524)
g25574(1) = AND(I24709, I24710)
g27085(1) = AND(g25835, g22494)
g28532(1) = AND(g27394, g20265)
g24707(1) = AND(g13295, g22997)
g25532(1) = NAND(g21360, g23363)
g25527(1) = NAND(g21294, g23462)
g22938(1) = AND(g19782, g19739)
g24706(1) = AND(g15910, g22996)
g23810(1) = NAND(I22973, I22974)
g23786(1) = NAND(I22945, I22946)
g25105(1) = AND(g13973, g23505)
g22681(1) = NAND(I21993, I21994)
g22663(1) = NAND(I21977, I21978)
g24624(1) = AND(g16524, g22867)
g26879(1) = OR(g25580, g25581)
g26878(1) = OR(g25578, g25579)
I24117(1) = OR(g23088, g23154, g23172)
I23755(1) = OR(g22904, g22927, g22980, g23444)
I26742(1) = OR(g23430, g23445, g23458, g23481)
I23756(1) = OR(g23457, g23480, g23494, g23511)
g26866(2) = OR(g20204, g20242, g24363)
g24916(1) = NAND(g19450, g23154)
g25779(2) = NAND(g19694, g24362)
g24942(1) = NAND(g20039, g23172)
g24917(1) = NAND(g19913, g23172)
g25018(1) = NAND(g20107, g23154)
g24918(1) = NAND(g136, g23088)
g24601(1) = NAND(g22957, g2965)
g24677(1) = NAND(g22957, g2975)
g24924(1) = NAND(g20007, g23172)
g24905(1) = NAND(g534, g23088)
g25002(1) = NAND(g19474, g23154)
g24621(1) = NAND(g22957, g2927)
I23961(2) = NAND(g23184, g13631)
I23585(2) = NAND(g22409, g4332)
g24972(1) = NAND(g19962, g23172)
g24950(1) = NAND(g19442, g23154)
g24906(1) = NAND(g8743, g23088)
g24383(1) = NOR(g22409, g22360)
g25425(1) = NAND(g20081, g23172)
g26256(2) = NOR(g23873, g25479)
g24631(2) = NOR(g20516, g20436, g20219, g22957)
I23949(2) = NAND(g23162, g13603)
g24933(1) = NAND(g19466, g23154)
g24567(1) = NAND(g22957, g2917)
g24662(1) = NAND(g22957, g2955)
I24461(2) = NAND(g23796, g14437)
I22923(1) = NAND(g21284, I22921)
I24363(2) = NAND(g23687, g14320)
g24932(1) = NAND(g19886, g23172)
g25540(1) = NOR(g22409, g22360)
g24925(1) = NAND(g20092, g23154)
I23978(2) = NAND(g23198, g13670)
I22922(1) = NAND(g14677, I22921)
g26212(2) = NOR(g23837, g25408)
I23985(2) = NAND(g22182, g482)
I23969(2) = NAND(g22202, g490)
I24383(2) = NAND(g23721, g14347)
g24988(1) = NAND(g546, g23088)
I23917(2) = NAND(g23975, g9333)
g25048(1) = NAND(g542, g23088)
I23600(2) = NAND(g22360, g4322)
I24438(2) = NAND(g23771, g14411)
I24414(2) = NAND(g23751, g14382)
g25019(1) = NAND(g20055, g23172)
g24570(1) = NAND(g22957, g2941)
g24576(1) = NAND(g22957, g2902)
g24951(1) = NAND(g199, g23088)
g25381(1) = NAND(g538, g23088)
g24943(1) = NAND(g20068, g23172)
g23683(1) = NOT(I22816)
g25167(1) = NOT(I24331)
g25259(1) = NOT(I24445)
g28041(1) = OR(g24145, g26878)
g28042(1) = OR(g24148, g26879)
g24168(1) = NOT(I23348)
g24178(1) = NOT(I23378)
g24174(1) = NOT(I23366)
g24181(1) = NOT(I23387)
g24172(1) = NOT(I23360)
g24161(1) = NOT(I23327)
g24177(1) = NOT(I23375)
g24171(1) = NOT(I23357)
g24163(1) = NOT(I23333)
g24170(1) = NOT(I23354)
g24185(1) = NOT(I23399)
g24164(1) = NOT(I23336)
g24173(1) = NOT(I23363)
g24162(1) = NOT(I23330)
g24179(1) = NOT(I23381)
g24180(1) = NOT(I23384)
g24175(1) = NOT(I23369)
g24183(1) = NOT(I23393)
g24166(1) = NOT(I23342)
g24176(1) = NOT(I23372)
g24184(1) = NOT(I23396)
g24169(1) = NOT(I23351)
g24182(1) = NOT(I23390)
g24165(1) = NOT(I23339)
g24167(1) = NOT(I23345)
g25751(1) = OR(g25061, g22098)
g29248(1) = OR(g28677, g18434)
g29223(1) = OR(g28341, g18131)
g24256(1) = OR(g22873, g18309)
g25728(1) = OR(g25076, g22011)
g25743(1) = OR(g25110, g22058)
g25599(1) = OR(g24914, g21721)
g29226(1) = OR(g28455, g18159)
g28076(1) = OR(g27098, g21878)
g25594(1) = OR(g24772, g21708)
g25741(1) = OR(g25178, g22056)
g25676(1) = OR(g24668, g21833)
g28070(1) = OR(g27050, g21867)
g25693(1) = OR(g24627, g18707)
g25661(1) = OR(g24754, g21786)
g25651(1) = OR(g24680, g21744)
g28077(1) = OR(g27120, g21879)
g25697(1) = OR(g25086, g21916)
g25650(1) = OR(g24663, g21743)
g25755(1) = OR(g25192, g22102)
g25595(1) = OR(g24835, g21717)
g26940(1) = OR(g25908, g21886)
g25709(1) = OR(g25014, g21960)
g25704(1) = OR(g25173, g21925)
g29230(1) = OR(g28107, g18202)
g25648(1) = OR(g24644, g21741)
g25731(1) = OR(g25128, g22014)
g28078(1) = OR(g27140, g21880)
g25739(1) = OR(g25149, g22054)
g25711(1) = OR(g25105, g21962)
g25703(1) = OR(g25087, g21922)
g25757(1) = OR(g25132, g22104)
g25729(1) = OR(g25091, g22012)
g25730(1) = OR(g25107, g22013)
g25679(1) = OR(g24728, g21836)
g29250(1) = OR(g28695, g18460)
g29275(1) = OR(g28165, g21868)
g25723(1) = OR(g25033, g22006)
g29235(1) = OR(g28110, g18260)
g25660(1) = OR(g24726, g21785)
g25726(1) = OR(g25148, g22009)
g25727(1) = OR(g25163, g22010)
g25677(1) = OR(g24684, g21834)
g25678(1) = OR(g24709, g21835)
g25671(1) = OR(g24637, g21828)
g25715(1) = OR(g25071, g21966)
g25674(1) = OR(g24755, g21831)
g25716(1) = OR(g25088, g21967)
g25675(1) = OR(g24769, g21832)
g25701(1) = OR(g25054, g21920)
g25713(1) = OR(g25147, g21964)
g29255(1) = OR(g28714, g18516)
g25732(1) = OR(g25201, g22017)
g25657(1) = OR(g24624, g21782)
g25746(1) = OR(g25217, g22063)
g25710(1) = OR(g25031, g21961)
g25591(1) = OR(g24642, g21705)
g25714(1) = OR(g25056, g21965)
g25680(1) = OR(g24794, g21839)
g25724(1) = OR(g25043, g22007)
g25718(1) = OR(g25187, g21971)
g25694(1) = OR(g24638, g18738)
g24240(1) = OR(g22861, g18251)
g25700(1) = OR(g25040, g21919)
g25691(1) = OR(g24536, g21890)
g28072(1) = OR(g27086, g21874)
g25712(1) = OR(g25126, g21963)
g25672(1) = OR(g24647, g21829)
g25695(1) = OR(g24998, g21914)
g29253(1) = OR(g28697, g18490)
g25758(1) = OR(g25151, g22105)
g29244(1) = OR(g28692, g18380)
g25645(1) = OR(g24679, g21738)
g29245(1) = OR(g28676, g18384)
g25658(1) = OR(g24635, g21783)
g28043(1) = OR(g27323, g21714)
g29251(1) = OR(g28679, g18464)
g25665(1) = OR(g24708, g21790)
g25592(1) = OR(g24672, g21706)
g25644(1) = OR(g24622, g21737)
g25662(1) = OR(g24656, g21787)
g25744(1) = OR(g25129, g22059)
g26938(1) = OR(g26186, g21883)
g25756(1) = OR(g25112, g22103)
g30334(1) = OR(g29837, g18143)
g25725(1) = OR(g25127, g22008)
g29228(1) = OR(g28426, g18173)
g25696(1) = OR(g25012, g21915)
g25685(1) = OR(g24476, g21866)
g29225(1) = OR(g28451, g18158)
g25760(1) = OR(g25238, g22109)
g24257(1) = OR(g22938, g18310)
g25673(1) = OR(g24727, g21830)
g25593(1) = OR(g24716, g21707)
g25752(1) = OR(g25079, g22099)
g29243(1) = OR(g28657, g18358)
g25740(1) = OR(g25164, g22055)
g29252(1) = OR(g28712, g18486)
g29227(1) = OR(g28456, g18169)
g25745(1) = OR(g25150, g22060)
g25753(1) = OR(g25165, g22100)
g25702(1) = OR(g25068, g21921)
g29240(1) = OR(g28655, g18328)
g25647(1) = OR(g24725, g21740)
g25699(1) = OR(g25125, g21918)
g29254(1) = OR(g28725, g18512)
g28074(1) = OR(g27119, g21876)
g29247(1) = OR(g28694, g18410)
g28071(1) = OR(g27085, g21873)
g25737(1) = OR(g25045, g22052)
g28075(1) = OR(g27083, g21877)
g25646(1) = OR(g24706, g21739)
g25597(1) = OR(g24892, g21719)
g29242(1) = OR(g28674, g18354)
g25659(1) = OR(g24707, g21784)
g25754(1) = OR(g25179, g22101)
g28073(1) = OR(g27097, g21875)
g24241(1) = OR(g22920, g18252)
g25698(1) = OR(g25104, g21917)
g26939(1) = OR(g25907, g21884)
g25596(1) = OR(g24865, g21718)
g25652(1) = OR(g24777, g21747)
g28053(1) = OR(g27393, g18168)
g29229(1) = OR(g28532, g18191)
g25649(1) = OR(g24654, g21742)
g25759(1) = OR(g25166, g22106)
g29241(1) = OR(g28638, g18332)
g25738(1) = OR(g25059, g22053)
g25664(1) = OR(g24681, g21789)
g26944(1) = OR(g26130, g18658)
g29246(1) = OR(g28710, g18406)
g25742(1) = OR(g25093, g22057)
g25643(1) = OR(g24602, g21736)
g25686(1) = OR(g24712, g21881)
g29249(1) = OR(g28658, g18438)
g25687(1) = OR(g24729, g21882)
g29256(1) = OR(g28597, g18533)
g28048(1) = OR(g27362, g18163)
g25717(1) = OR(g25106, g21968)
g25598(1) = OR(g24904, g21720)
g25666(1) = OR(g24788, g21793)
g25663(1) = OR(g24666, g21788)
g25027(2) = NOT(I24191)
g27907(16) = OR(g17424, g26770)
I24237(1) = NOT(g23823)
g25249(1) = NOT(g22228)
g25248(1) = NOT(g22228)
g25552(1) = NOT(g22594)
g27084(1) = NOT(g26673)
g27800(16) = OR(g17321, g26703)
g25786(1) = NOT(g24518)
I28576(1) = NOT(g28431)
g24431(1) = NOT(g22722)
g24920(1) = NOT(I24089)
g25380(1) = NOT(g23776)
g29744(1) = NOT(g28431)
g25206(1) = NOT(g23613)
g27511(3) = NOR(g22137, g26866, g20277)
g25513(1) = NOT(g23870)
g25505(1) = NOT(g22228)
I27192(1) = NOT(g27662)
g25369(1) = NOT(g22228)
g25424(1) = NOT(g23800)
g27008(1) = OR(g26866, g21370, I25736)
g25641(1) = NOT(I24784)
g29507(1) = NOT(g28353)
g27983(1) = NOT(g26725)
g27837(16) = OR(g17401, g26725)
g24417(1) = NOT(g22171)
g25548(1) = NOT(g22550)
I25586(1) = NOT(g25537)
g24836(2) = NOT(I24008)
g25533(1) = NOT(g22550)
g25298(1) = NOT(g23760)
g27779(16) = OR(g17317, g26694)
g25232(1) = NOT(g22228)
I26004(1) = NOT(g26818)
g25198(1) = NOT(g22228)
g25528(1) = NOT(g22594)
g25250(4) = NOT(I24434)
g23453(2) = NOT(I22576)
g27091(1) = NOT(g26725)
g25171(1) = NOT(g22228)
g25886(1) = NOT(g24537)
g27858(16) = OR(g17405, g26737)
g30322(2) = NOT(g28431)
I25327(1) = NOT(g24641)
g25322(1) = NOT(I24497)
g25158(1) = NOT(g22228)
g27742(16) = OR(g17292, g26673)
g25561(1) = NOT(g22550)
g25241(1) = NOT(g23651)
g25260(1) = NOT(I24448)
g25272(1) = NOT(g23715)
I25594(1) = NOT(g25531)
g24759(1) = NOT(g23003)
g25289(1) = NOT(g22228)
g24891(1) = NOT(g23231)
g25288(1) = NOT(g22228)
g26424(58) = NOT(I25356)
g25525(1) = NOT(g22550)
g25558(1) = NOT(g22594)
g25830(1) = NOT(g24485)
g25893(1) = NOT(g24541)
g25544(1) = NOT(g22594)
g24869(2) = NOT(I24041)
g24483(1) = NOT(I23688)
g25296(1) = NOT(g23745)
g25267(1) = NOT(g22228)
g25064(2) = NOT(I24228)
g24866(2) = NOT(I24038)
g24452(1) = NOT(g22722)
g28121(2) = NOT(g27093)
g25689(1) = OR(g24849, g21888)
g29707(1) = NOT(g28504)
g25266(1) = NOT(g22228)
g27886(16) = OR(g14438, g26759)
g25524(1) = NOT(g22228)
g24405(1) = NOT(g22722)
g25642(1) = NOT(I24787)
g31243(1) = NOT(g29933)
g27971(1) = NOT(g26673)
g29597(1) = NOT(g28444)
g25560(1) = NOT(g22550)
g26187(2) = NOT(I25190)
g25917(3) = OR(g22524, g24518)
g24489(1) = NOT(I23694)
g25555(1) = NOT(g22550)
g27112(1) = NOT(g26793)
g24356(1) = NOT(g22594)
g25185(1) = NOT(g22228)
g25284(1) = NOT(I24474)
I26654(1) = NOT(g27576)
g25566(1) = NOT(g22550)
g25180(1) = NOT(g23529)
I25359(1) = NOT(g24715)
g24368(1) = NOT(g22228)
g24850(2) = NOT(I24022)
g27989(1) = NOT(g26759)
g25554(1) = NOT(g22550)
I24281(1) = NOT(g23440)
g24379(1) = NOT(g22550)
g24386(1) = NOT(g22594)
g24429(1) = NOT(g22722)
g24428(1) = NOT(g22722)
g25214(1) = NOT(g22228)
g28127(2) = NOT(g27102)
g25538(1) = NOT(g22594)
g27994(1) = NOT(g26793)
I24278(1) = NOT(g23440)
g25849(1) = NOT(g24491)
g24365(1) = NOT(g22594)
g25221(1) = NOT(g23653)
g27976(1) = NOT(g26703)
g24375(1) = NOT(g22722)
g24425(1) = NOT(g22722)
g24911(1) = NOT(I24078)
g25325(1) = NOT(g22228)
g24477(1) = NOT(I23680)
g27937(16) = OR(g14506, g26793)
g25506(1) = NOT(g22228)
g24364(1) = NOT(g22722)
g25265(1) = NOT(I24455)
g25168(1) = NOT(I24334)
g25240(1) = NOT(g23650)
g27984(1) = NOT(g26737)
I26667(1) = NOT(g27585)
g25563(1) = NOT(g22594)
g24424(1) = NOT(g22722)
g24893(2) = NOT(I24060)
g25324(1) = NOT(g22228)
g27101(1) = NOT(g26770)
g25140(1) = NOT(g22228)
g25911(3) = OR(g22514, g24510)
g25451(1) = NOT(g22228)
g25690(1) = OR(g24864, g21889)
g27092(1) = NOT(g26737)
g25370(1) = NOT(g22228)
g24419(1) = NOT(g22722)
g24418(1) = NOT(g22722)
g25688(1) = OR(g24812, g21887)
g24466(1) = NOT(I23671)
g24229(1) = AND(g896, g22594)
g25547(1) = NOT(g22550)
g25481(1) = NOT(g22228)
g25297(1) = NOT(g23746)
g25640(1) = NOT(I24781)
g25546(1) = NOT(g22550)
I28128(1) = NOT(g28314)
g24438(1) = NOT(g22722)
g27100(1) = NOT(g26759)
g27599(1) = AND(g26337, g20033)
g29343(1) = NOT(g28174)
g31509(3) = NAND(g599, g29933, g12323)
g25231(1) = NOT(g22228)
g24407(1) = NOT(g22594)
g23684(1) = NOT(I22819)
g25480(1) = NOT(g22228)
g25287(1) = NOT(g22228)
g28508(1) = NOT(I26989)
g25286(1) = NOT(g22228)
g27990(1) = NOT(g26770)
g25410(1) = NOT(g22228)
g24359(1) = NOT(g22550)
g24358(1) = NOT(g22550)
g25465(1) = NOT(g23824)
g25517(1) = NOT(g22228)
g25523(1) = NOT(g22550)
g24360(1) = NOT(g22228)
g25781(1) = NOT(g24510)
g24367(1) = NOT(g22550)
g24394(1) = NOT(g22228)
g27089(1) = NOT(g26703)
g27088(1) = NOT(g26694)
g29916(3) = NOR(g8681, g28504, g11083)
g24377(1) = NOT(g22594)
g25409(1) = NOT(g22228)
g24366(1) = NOT(g22594)
g24481(1) = NOT(I23684)
g24298(1) = AND(g4392, g22550)
g24490(1) = NOT(g22594)
g26326(1) = NOT(g24872)
g24376(1) = NOT(g22722)
g29778(3) = NAND(g294, g28444, g23204)
g24426(1) = NOT(g22722)
g25553(1) = NOT(g22550)
g25326(1) = NOT(g22228)
g29333(1) = NOT(g28167)
g29679(3) = NAND(g153, g28353, g23042)
g25452(1) = NOT(g22228)
g24819(1) = NOT(I23998)
g25051(2) = NOT(I24215)
g27975(1) = NOT(g26694)
g26865(1) = NOR(g25328, g25290)
g24314(1) = AND(g4515, g22228)
g24287(1) = AND(g4401, g22550)
g24307(1) = AND(g4486, g22228)
g25357(8) = AND(g23810, g23786)
g30149(1) = AND(g28605, g21248)
g24286(1) = AND(g4405, g22550)
g24306(1) = AND(g4483, g22228)
g30133(1) = AND(g28591, g21179)
g28208(1) = OR(g27025, g27028)
g24187(1) = AND(g305, g22722)
g27265(1) = AND(g26785, g26759)
g26800(1) = OR(g24922, g24929)
g30112(1) = AND(g28566, g20919)
g26857(1) = AND(g25062, g25049)
g24217(1) = AND(g18200, g22594)
g30096(1) = AND(g28546, g20770)
g28616(1) = AND(g27532, g20551)
g28313(1) = AND(g27231, g19766)
g27615(1) = AND(g26789, g26770)
g24223(1) = AND(g239, g22594)
g24321(1) = AND(g4558, g22228)
g23778(1) = NAND(I22922, I22923)
g31144(1) = OR(g29477, g28193)
g24186(1) = AND(g18102, g22722)
g25765(1) = AND(g24989, g24973)
g24688(9) = AND(g22681, g22663)
g27600(1) = AND(g26755, g26725)
g28185(1) = AND(g27026, g19435)
g30579(1) = OR(g30173, g14571)
g24230(1) = AND(g901, g22594)
g24293(1) = AND(g4438, g22550)
g30145(1) = AND(g28603, g21247)
g27614(1) = AND(g26785, g26759)
g29324(1) = AND(g29078, g18883)
g30161(1) = AND(g28614, g21275)
g28415(1) = AND(g27250, g19963)
g24193(1) = AND(g336, g22722)
g24222(1) = AND(g262, g22594)
g28211(1) = OR(g27029, g27034)
g30078(1) = AND(g28526, g20667)
g30086(1) = AND(g28536, g20704)
g30125(1) = AND(g28581, g21056)
g29367(1) = AND(g8575, g28325)
g30158(1) = AND(g28613, g21274)
g26293(1) = OR(g24550, g24555)
g27252(1) = AND(g26733, g26703)
g26305(1) = OR(g24556, g24564)
g24320(1) = AND(g6973, g22228)
g24952(1) = OR(g21326, g21340, I24117)
g25769(1) = NOR(g25453, g25414)
g28132(1) = OR(g27932, g27957)
g27634(1) = AND(g26805, g26793)
g24292(1) = AND(g4443, g22550)
g24327(1) = AND(g4549, g22228)
g24283(1) = AND(g4411, g22550)
g24303(1) = AND(g4369, g22228)
g29376(1) = AND(g14002, g28504)
g25778(1) = NOR(g25459, g25420)
g24192(1) = AND(g311, g22722)
g30124(1) = AND(g28580, g21055)
g24326(1) = AND(g4552, g22228)
g25985(1) = NAND(g24631, g23956)
g28216(1) = OR(g27036, g27043)
g30075(1) = AND(g28525, g20662)
g24311(1) = AND(g4498, g22228)
g30118(1) = AND(g28574, g21050)
g30101(1) = AND(g28551, g20780)
g30064(1) = AND(g28517, g20630)
g26485(1) = AND(g24968, g10502)
g24302(1) = AND(g15124, g22228)
g28440(1) = AND(g27274, g20059)
g26574(1) = NOR(g24887, g24861)
g30935(1) = AND(g8808, g29745)
g25784(1) = NOR(g25507, g25485)
g24331(1) = AND(g6977, g22228)
g30083(1) = AND(g28533, g20698)
g26852(1) = AND(g24975, g24958)
g30139(1) = AND(g28596, g21184)
g30138(1) = AND(g28595, g21182)
g26546(1) = NOR(g24858, g24846)
g26573(1) = NOR(g24897, g24884)
g26484(1) = AND(g24946, g8841)
g25785(1) = NOR(g25488, g25462)
g26809(1) = OR(g24930, g24939)
g31654(1) = AND(g29325, g13062)
g29937(1) = AND(g13044, g29196)
g24228(1) = AND(g862, g22594)
g29363(1) = AND(g8458, g28444)
g26781(1) = OR(g24913, g24921)
g28301(1) = AND(g27224, g19750)
g24310(1) = AND(g4495, g22228)
g25800(1) = NOR(g25518, g25510)
g28427(1) = AND(g27258, g20008)
g27259(1) = AND(g26755, g26725)
g24317(1) = AND(g4534, g22228)
g24323(1) = AND(g4546, g22228)
g24299(1) = AND(g4456, g22550)
g26398(1) = AND(g24946, g10474)
g30107(1) = AND(g28560, g20909)
g27598(1) = AND(g25899, g10475)
g24316(1) = AND(g4527, g22228)
g30135(1) = AND(g28592, g21180)
g26613(1) = AND(g1361, g24518)
g30049(1) = AND(g13114, g28167)
g29746(1) = AND(g28279, g20037)
g24199(1) = AND(g355, g22722)
g24198(1) = AND(g351, g22722)
g24330(1) = AND(g18661, g22228)
g26603(1) = NOR(g24908, g24900)
g26515(1) = NOR(g24843, g24822)
g26025(1) = NAND(g22405, g24631)
g24225(1) = AND(g246, g22594)
g27260(1) = AND(g26766, g26737)
g30121(1) = AND(g28577, g21052)
g25774(1) = OR(g25223, g12043)
g29834(1) = AND(g28368, g23278)
g27270(1) = AND(g26805, g26793)
g24322(1) = AND(g4423, g22228)
g24295(1) = AND(g4434, g22550)
g24289(1) = AND(g4427, g22550)
g24309(1) = AND(g4480, g22228)
g24288(1) = AND(g4417, g22550)
g27595(1) = AND(g26733, g26703)
g24224(1) = AND(g269, g22594)
g24308(1) = AND(g4489, g22228)
g31252(1) = AND(g29643, g20101)
g26861(1) = AND(g25021, g25003)
g27266(1) = AND(g26789, g26770)
g28135(1) = OR(g27959, g27963)
g27588(1) = AND(g26690, g26673)
g30099(1) = AND(g28549, g20776)
g24195(1) = AND(g74, g22722)
g30098(1) = AND(g28548, g20774)
g26871(1) = AND(g25038, g25020)
g24189(1) = AND(g324, g22722)
g24188(1) = AND(g316, g22722)
g24294(1) = AND(g4452, g22550)
g26872(1) = NOR(g25411, g25371)
g24219(1) = AND(g225, g22594)
g24218(1) = AND(g872, g22594)
g30151(1) = AND(g28607, g21249)
g30172(1) = AND(g28625, g21286)
g27594(1) = AND(g26721, g26694)
g28178(1) = AND(g27019, g19397)
g24194(1) = AND(g106, g22722)
g30120(1) = AND(g28576, g21051)
g24313(1) = AND(g4504, g22228)
g24285(1) = AND(g4388, g22550)
g24305(1) = AND(g4477, g22228)
g28442(1) = AND(g27278, g20072)
g30095(1) = AND(g28545, g20768)
g30671(1) = AND(g29319, g22317)
g29508(1) = OR(g28152, g27041)
g26873(1) = NOR(g25374, g25331)
g30089(1) = AND(g28538, g20709)
g28134(1) = OR(g27958, g27962)
g30126(1) = AND(g28582, g21058)
g29513(1) = AND(g28448, g14095)
g24284(1) = AND(g4375, g22550)
g24304(1) = AND(g12875, g22228)
g25770(1) = NOR(g25417, g25377)
g24333(1) = AND(g4512, g22228)
g30111(1) = AND(g28565, g20917)
g30094(1) = AND(g28544, g20767)
g24312(1) = AND(g4501, g22228)
g29378(1) = AND(g28137, g22493)
g24329(1) = AND(g4462, g22228)
g30066(1) = AND(g28518, g20636)
g24328(1) = AND(g4567, g22228)
g29706(1) = OR(g28198, g27208)
g25767(1) = OR(g25207, g12015)
g26278(1) = OR(g24545, g24549)
g29359(1) = NOR(g7528, g28167)
g30131(1) = AND(g28589, g21178)
g29793(1) = OR(g28237, g27247)
g25777(1) = NOR(g25482, g25456)
g28183(1) = AND(g27024, g19421)
g29924(1) = AND(g13031, g29190)
g24332(1) = AND(g4459, g22228)
g29330(1) = AND(g29114, g18894)
g27648(1) = AND(g25882, g8974)
g24221(1) = AND(g232, g22594)
g26751(1) = OR(g24903, g24912)
g29375(1) = AND(g13946, g28370)
g30084(1) = AND(g28534, g20700)
g30110(1) = AND(g28564, g20916)
g27612(1) = AND(g25887, g8844)
g27251(1) = AND(g26721, g26694)
g24325(1) = AND(g4543, g22228)
g26813(1) = OR(g24940, g24949)
g24291(1) = AND(g18660, g22550)
g27246(1) = AND(g26690, g26673)
g25772(1) = AND(g24944, g24934)
g24191(1) = AND(g319, g22722)
g29668(1) = AND(g28527, g14255)
g24324(1) = AND(g4540, g22228)
g26863(1) = AND(g24974, g24957)
g28138(1) = OR(g27964, g27968)
g26516(1) = AND(g24968, g8876)
g30287(1) = OR(g28653, g27677)
g24220(1) = AND(g255, g22594)
g30137(1) = AND(g28594, g21181)
g29494(1) = AND(g9073, g28479)
g30291(1) = OR(g28672, g27685)
g30122(1) = AND(g28578, g21054)
g24319(1) = AND(g4561, g22228)
g24318(1) = AND(g4555, g22228)
g24227(1) = AND(g890, g22594)
g28626(1) = AND(g27542, g20573)
g29583(1) = OR(g28182, g27099)
g24301(1) = AND(g6961, g22228)
g26606(1) = AND(g1018, g24510)
g24290(1) = AND(g4430, g22550)
g30109(1) = AND(g28562, g20912)
g30108(1) = AND(g28561, g20910)
g28212(1) = OR(g27030, g27035)
g30982(1) = AND(g8895, g29933)
g24226(1) = AND(g446, g22594)
g29570(1) = AND(g2763, g28598)
g24297(1) = AND(g4455, g22550)
g24190(1) = AND(g329, g22722)
g30062(1) = AND(g13129, g28174)
g28171(1) = AND(g27016, g19385)
g24296(1) = AND(g4382, g22550)
g24197(1) = AND(g347, g22722)
g30051(1) = AND(g28513, g20604)
g26545(1) = NOR(g24881, g24855)
g24315(1) = AND(g4521, g22228)
g29361(1) = NOR(g7553, g28174)
g25780(1) = AND(g25532, g25527)
g24196(1) = AND(g333, g22722)
g29329(1) = AND(g7995, g28353)
g27601(1) = AND(g26766, g26737)
g24300(1) = AND(g15123, g22228)
g26052(1) = NAND(g22714, g24662, g22921)
g25974(1) = NAND(g24576, g22837)
g25856(8) = OR(g25518, g25510, g25488, g25462)
g25504(1) = NOR(g22550, g7222)
g25141(1) = NOR(g22228, g10334)
g26657(8) = OR(g24908, g24900, g24887, g24861)
g24561(2) = OR(I23755, I23756)
g25953(1) = NAND(g22756, g24570, g22688)
g26616(8) = OR(g24881, g24855, g24843, g24822)
I25612(1) = OR(g25567, g25568, g25569, g25570)
I25613(1) = OR(g25571, g25572, g25573, g25574)
g26636(8) = OR(g24897, g24884, g24858, g24846)
g25996(1) = NAND(g24601, g22838)
g26053(1) = NAND(g22875, g24677, g22941)
g25805(8) = OR(g25453, g25414, g25374, g25331)
g25995(1) = NAND(g24621, g22853)
g25984(1) = NAND(g24567, g22668)
g25839(8) = OR(g25507, g25485, g25459, g25420)
g25791(8) = OR(g25411, g25371, g25328, g25290)
g25821(8) = OR(g25482, g25456, g25417, g25377)
I25242(2) = NAND(g490, g24744)
I23979(1) = NAND(g23198, I23978)
I23980(1) = NAND(g13670, I23978)
I23963(1) = NAND(g13631, I23961)
I25219(2) = NAND(g482, g24718)
I24462(1) = NAND(g23796, I24461)
I24463(1) = NAND(g14437, I24461)
I24364(1) = NAND(g23687, I24363)
I24365(1) = NAND(g14320, I24363)
I24439(1) = NAND(g23771, I24438)
I24440(1) = NAND(g14411, I24438)
I25907(2) = NAND(g26256, g24782)
I23962(1) = NAND(g23184, I23961)
I23951(1) = NAND(g13603, I23949)
g29660(1) = NAND(g28448, g9582)
I23950(1) = NAND(g23162, I23949)
I23601(1) = NAND(g22360, I23600)
I23602(1) = NAND(g4322, I23600)
I24384(1) = NAND(g23721, I24383)
I24385(1) = NAND(g14347, I24383)
I23586(1) = NAND(g22409, I23585)
I23587(1) = NAND(g4332, I23585)
I23970(1) = NAND(g22202, I23969)
I23971(1) = NAND(g490, I23969)
I25845(2) = NAND(g26212, g24799)
I23987(1) = NAND(g482, I23985)
I23986(1) = NAND(g22182, I23985)
I24415(1) = NAND(g23751, I24414)
I23918(1) = NAND(g23975, I23917)
I23919(1) = NAND(g9333, I23917)
I24416(1) = NAND(g14382, I24414)
g25114(1) = NOT(I24278)
g30381(1) = OR(g30126, g18497)
g30360(1) = OR(g30145, g18386)
g30384(1) = OR(g30101, g18517)
g30348(1) = OR(g30083, g18329)
g29236(1) = OR(g28313, g18287)
g30335(1) = OR(g29746, g18174)
g29239(1) = OR(g28427, g18297)
g29279(1) = OR(g28442, g18741)
g30370(1) = OR(g30135, g18440)
g30366(1) = OR(g30122, g18417)
g30336(1) = OR(g29324, g18203)
g30369(1) = OR(g30066, g18439)
g29276(1) = OR(g28616, g18709)
g31894(1) = OR(g30671, g21870)
g29237(1) = OR(g28185, g18289)
g30378(1) = OR(g30125, g18487)
g29278(1) = OR(g28626, g18740)
g30350(1) = OR(g30118, g18334)
g30383(1) = OR(g30138, g18513)
g30377(1) = OR(g30124, g18472)
g30362(1) = OR(g30120, g18392)
g30456(1) = OR(g29378, g21869)
g30371(1) = OR(g30099, g18445)
g30368(1) = OR(g30098, g18435)
g30375(1) = OR(g30149, g18466)
g30349(1) = OR(g30051, g18333)
g29238(1) = OR(g28178, g18292)
g30379(1) = OR(g30089, g18491)
g30382(1) = OR(g30137, g18498)
g30363(1) = OR(g30121, g18407)
g30356(1) = OR(g30096, g18365)
g30365(1) = OR(g30158, g18412)
g29232(1) = OR(g28183, g18231)
g30374(1) = OR(g30078, g18465)
g30342(1) = OR(g29330, g18261)
g30364(1) = OR(g30086, g18411)
g30353(1) = OR(g30095, g18355)
g30372(1) = OR(g30110, g18446)
g30354(1) = OR(g30064, g18359)
g30333(1) = OR(g29834, g21699)
g30387(1) = OR(g30151, g18524)
g30357(1) = OR(g30107, g18366)
g30358(1) = OR(g30108, g18381)
g30367(1) = OR(g30133, g18418)
g30359(1) = OR(g30075, g18385)
g30351(1) = OR(g30084, g18339)
g31866(1) = OR(g31252, g18142)
g30373(1) = OR(g30111, g18461)
g30355(1) = OR(g30131, g18360)
g30386(1) = OR(g30139, g18523)
g29233(1) = OR(g28171, g18234)
g30376(1) = OR(g30112, g18471)
g29234(1) = OR(g28415, g18239)
g30385(1) = OR(g30172, g18518)
g30361(1) = OR(g30109, g18391)
g29231(1) = OR(g28301, g18229)
g30380(1) = OR(g30161, g18492)
g30352(1) = OR(g30094, g18340)
g29277(1) = OR(g28440, g18710)
g28713(1) = NOT(g27907)
g29134(6) = NAND(g9762, g27907)
g28678(1) = NOT(g27800)
I25105(1) = NOT(g25284)
I25161(1) = NOT(g24920)
g26811(1) = NOT(g25206)
I27492(1) = NOT(g27511)
g29118(2) = NAND(g27886, g9755)
I25576(1) = NOT(g25296)
g26365(11) = OR(g25504, g25141)
I24759(1) = NOT(g24229)
I25598(1) = NOT(g25424)
g28709(1) = NOT(I27192)
g28830(2) = NAND(g27886, g7451, g7369)
g28119(1) = NOT(g27008)
I25680(1) = NOT(g25641)
I25391(1) = NOT(g24483)
g28824(2) = NAND(g27779, g7356, g1772)
g26260(1) = NOT(g24759)
g28693(1) = NOT(g27837)
g28765(2) = NAND(g27800, g7374, g7280)
g26856(1) = NOT(I25586)
g26831(1) = NOT(g24836)
g28861(2) = NAND(g27837, g7405, g1906)
g28675(1) = NOT(g27779)
g28942(2) = NAND(g27858, g2331, g7335)
I25567(1) = NOT(g25272)
g27320(2) = NOT(I26004)
g29045(1) = NOT(g27779)
g29121(6) = NAND(g9755, g27886)
g29060(6) = NAND(g9649, g27800)
g25869(1) = NOT(g25250)
g29157(6) = NAND(g9835, g27937)
g31227(1) = NOT(g29744)
I24396(1) = NOT(g23453)
g28780(2) = NAND(g27742, g7308, g1636)
g25242(1) = NOT(g23684)
g29097(6) = NAND(g9700, g27858)
g28896(2) = NAND(g27837, g1936, g1862)
g29151(1) = NOT(g27858)
g28962(2) = NAND(g27886, g2040, g7369)
g26364(1) = NOT(I25327)
g29085(6) = NAND(g9694, g27837)
g25783(1) = NOT(g25250)
g29044(1) = NOT(g27742)
I25555(1) = NOT(g25241)
g26816(1) = NOT(g25260)
I25366(1) = NOT(g24477)
I25779(1) = NOT(g26424)
g29049(6) = NAND(g9640, g27779)
g28180(1) = OR(g20242, g27511)
g28935(2) = NAND(g27800, g2227, g7328)
g26837(1) = NOT(g24869)
g27660(1) = AND(g24688, g26424, g22763)
I25115(1) = NOT(g25322)
I24393(1) = NOT(g23453)
g25837(1) = NOT(g25064)
g26836(1) = NOT(g24866)
I25692(1) = NOT(g25689)
g28927(2) = NAND(g27837, g1906, g7322)
I25005(1) = NOT(g24417)
g29001(2) = NAND(g27937, g2599, g7431)
g28843(2) = NAND(g27907, g7456, g7387)
g29150(1) = NOT(g27886)
I25683(1) = NOT(g25642)
g28874(2) = NAND(g27907, g7424, g2421)
g31134(3) = NOR(g8033, g29679, g24732)
I26406(1) = NOT(g26187)
I25689(1) = NOT(g25688)
I25380(1) = NOT(g24481)
g29046(2) = NAND(g27779, g9640)
g27011(1) = NOT(g25917)
I25677(1) = NOT(g25640)
I25399(1) = NOT(g24489)
g27730(1) = NOT(g26424)
g28867(2) = NAND(g27800, g2227, g2153)
g29018(6) = NAND(g9586, g27742)
g28903(2) = NAND(g27800, g2197, g7280)
g25073(2) = NOT(I24237)
g28147(1) = NOT(I26654)
g26718(1) = NOT(g25168)
I25541(1) = NOT(g25180)
g31262(3) = NAND(g767, g29916, g11679)
g29169(1) = NOT(g27886)
I25351(1) = NOT(g24466)
g25115(1) = NOT(I24281)
g27108(3) = OR(g22522, g25911)
g28837(2) = NAND(g27800, g7374, g2197)
g28907(2) = NAND(g27858, g2361, g2287)
I24839(1) = NOT(g24298)
g29131(2) = NAND(g27907, g9762)
g29117(1) = NOT(g27886)
I24920(1) = NOT(g25513)
g29014(1) = NOT(g27742)
g27122(3) = OR(g22537, g25917)
g29116(1) = NOT(g27837)
g28977(2) = NAND(g27937, g2629, g2555)
I25591(1) = NOT(g25380)
g29130(1) = NOT(g27907)
g30325(1) = NOT(I28576)
I25146(1) = NOT(g24911)
I25562(1) = NOT(g25250)
g28840(2) = NAND(g27858, g7380, g2287)
g28783(2) = NAND(g27779, g7315, g1728)
g29153(1) = NOT(g27937)
I25095(1) = NOT(g25265)
g26832(1) = NOT(g24850)
g28156(1) = NOT(I26667)
I26936(1) = NOT(g27599)
I26710(1) = NOT(g27511)
g28853(2) = NAND(g27742, g1636, g7252)
I25786(1) = NOT(g26424)
I28913(1) = NOT(g30322)
g27009(1) = NOT(g25911)
I25790(1) = NOT(g26424)
I25695(1) = NOT(g25690)
g28827(2) = NAND(g27837, g7362, g1862)
g29152(1) = NOT(g27907)
g28914(2) = NAND(g27937, g7462, g2555)
g28871(2) = NAND(g27858, g7418, g2331)
g26824(1) = NOT(g25298)
g28758(2) = NAND(g27779, g7356, g7275)
g26860(1) = NOT(I25594)
g29081(1) = NOT(g27837)
g29094(2) = NAND(g27858, g9700)
g28973(2) = NAND(g27907, g2465, g7387)
g28966(2) = NAND(g27858, g2361, g7380)
I25606(1) = NOT(g25465)
g29897(1) = NOT(I28128)
g28892(2) = NAND(g27779, g1772, g7275)
g29149(1) = NOT(g27837)
g28726(1) = NOT(g27937)
g28987(2) = NAND(g27886, g2070, g7411)
g28820(2) = NAND(g27742, g1668, g1592)
g28911(2) = NAND(g27907, g7456, g2465)
g29057(2) = NAND(g27800, g9649)
g28711(1) = NOT(g27886)
g32201(1) = NOT(g31509)
I25579(1) = NOT(g25297)
g29129(1) = NOT(g27858)
g29128(1) = NOT(g27800)
g29082(2) = NAND(g27837, g9694)
g28955(2) = NAND(g27837, g1936, g7362)
g32296(3) = NOR(g9044, g31509, g12259)
g29056(1) = NOT(g27800)
g29080(1) = NOT(g27779)
g25838(1) = NOT(g25250)
g28796(2) = NAND(g27858, g7418, g7335)
g28885(2) = NAND(g27742, g1668, g7268)
I26409(1) = NOT(g26187)
g28950(2) = NAND(g27937, g7490, g2599)
g29171(1) = NOT(g27937)
g28946(2) = NAND(g27907, g2495, g2421)
g29079(1) = NOT(g27742)
g31233(3) = NOR(g8522, g29778, g24825)
g28920(2) = NAND(g27779, g1802, g7315)
g26814(1) = NOT(g25221)
g26841(1) = NOT(g24893)
I25369(1) = NOT(g24891)
g28755(2) = NAND(g27742, g7268, g1592)
g28857(2) = NAND(g27779, g1802, g1728)
g29093(1) = NOT(g27858)
g29015(2) = NAND(g27742, g9586)
I25552(1) = NOT(g25240)
g28994(2) = NAND(g27907, g2495, g7424)
g25790(1) = NOT(g25027)
g29170(1) = NOT(g27907)
g28736(2) = NAND(g27742, g7308, g7252)
g31239(1) = NOT(g29916)
g29177(1) = NOT(g27937)
g28786(2) = NAND(g27837, g7405, g7322)
g26483(1) = NOT(I25359)
g28696(1) = NOT(g27858)
g31138(1) = NOT(g29778)
g28900(2) = NAND(g27886, g7451, g2040)
g29092(1) = NOT(g27800)
g29025(2) = NAND(g27937, g2629, g7462)
g28793(2) = NAND(g27800, g7328, g2153)
g31013(1) = NOT(g29679)
g28931(2) = NAND(g27886, g2070, g1996)
g28656(1) = NOT(g27742)
g28877(2) = NAND(g27937, g7490, g7431)
g29115(1) = NOT(g27779)
g28864(2) = NAND(g27886, g7411, g1996)
g25820(1) = NOT(g25051)
g26827(1) = NOT(g24819)
g29154(2) = NAND(g27937, g9835)
g27703(1) = NOR(g9607, g25791)
g24798(1) = NAND(I23962, I23963)
I26960(1) = AND(g24995, g26424, g22698)
g27010(1) = NOR(g6052, g25839)
g26356(1) = AND(g15581, g25523)
g28149(1) = NOR(g27598, g27612)
g27666(1) = AND(g26865, g23521)
g26380(1) = AND(g19572, g25547)
g27969(1) = NOR(g7170, g25821)
g26236(4) = AND(g25357, g6856, g7586, g7558)
g26651(1) = AND(g22707, g24425)
g26513(1) = AND(g19501, g24365)
I27409(1) = AND(g25556, g26424, g22698)
g28255(1) = AND(g8515, g27983)
g27368(1) = NOR(g8119, g26657)
g26195(4) = AND(g25357, g6856, g11709, g7558)
g26148(4) = AND(g25357, g11724, g11709, g11686)
g27768(1) = NOR(g9264, g25805)
g26218(4) = AND(g25357, g6856, g7586, g11686)
g25199(1) = NAND(I24364, I24365)
I27381(1) = AND(g25549, g26424, g22698)
g27499(1) = NOR(g9095, g26636)
g26993(1) = NOR(g5360, g25805)
g27973(1) = NOR(g7187, g25839)
g31020(1) = OR(g29375, g28164)
g29613(1) = AND(g28208, g19763)
g26379(1) = AND(g19904, g25546)
g26378(1) = AND(g19576, g25544)
g27992(1) = AND(g26800, g23964)
g28524(1) = AND(g6821, g27084)
g27966(1) = NOR(g7153, g25805)
g27261(1) = OR(g24544, g25996)
g27241(1) = OR(g24584, g25984)
g30730(1) = AND(g26346, g29778)
g27960(1) = NOR(g7134, g25791)
g31474(1) = OR(g29668, g13583)
g25096(1) = AND(g23778, g20560)
g32197(1) = AND(g31144, g20088)
g26976(1) = NOR(g5016, g25791)
g26261(2) = AND(g24688, g10678, g8778, g8757)
g28567(1) = AND(g6832, g27101)
g32019(1) = AND(g30579, g22358)
g27587(1) = NAND(g24917, g25018, g24918, g26857)
g26753(1) = AND(g16024, g24452)
g26213(4) = AND(g25357, g11724, g7586, g7558)
g30080(1) = AND(g28121, g20674)
g26650(1) = AND(g10796, g24424)
g26393(1) = AND(g19467, g25558)
g28284(1) = AND(g11398, g27994)
g25258(1) = NAND(I24439, I24440)
g26281(2) = AND(g24688, g8812, g8778, g8757)
g26259(1) = AND(g24430, g25232)
g26258(1) = AND(g12875, g25231)
g27337(1) = NOR(g8334, g26616)
g27875(1) = NOR(g9875, g25821)
g26244(2) = AND(g24688, g8812, g10658, g8757)
g26171(4) = AND(g25357, g6856, g11709, g11686)
g27063(1) = NOR(g26485, g26516)
I26972(1) = AND(g25011, g26424, g22698)
g26226(2) = AND(g24688, g8812, g10658, g10627)
g26166(4) = AND(g25357, g11724, g11709, g7558)
g27828(1) = NOR(g9892, g25856)
g27652(1) = NOR(g3355, g26636)
g27253(1) = OR(g24661, g26052)
g27364(1) = NOR(g8426, g26616)
g27354(1) = NOR(g8064, g26636)
g29629(1) = AND(g28211, g19779)
g27924(1) = NOR(g9946, g25839)
g30918(1) = AND(g8681, g29707)
g26295(1) = AND(g13070, g25266)
g27731(1) = NOR(g9229, g25791)
g26336(1) = AND(g10307, g25480)
g27553(1) = AND(g26293, g23353)
g24807(1) = NAND(I23979, I23980)
g27564(1) = AND(g26305, g23378)
g25236(1) = NAND(I24415, I24416)
g26571(1) = AND(g10472, g24386)
g26308(1) = AND(g6961, g25289)
g27673(1) = AND(g25769, g23541)
g31014(1) = OR(g29367, g28160)
g29377(1) = AND(g28132, g19387)
g30023(1) = AND(g28508, g20570)
I27429(1) = AND(g25562, g26424, g22698)
g27613(1) = NAND(g24942, g24933, g25048, g26871)
g26610(1) = AND(g14198, g24405)
g27691(1) = AND(g25778, g23609)
g31527(1) = AND(g7553, g29343)
g27927(1) = NOR(g9621, g25856)
g27877(1) = NOR(g9397, g25839)
g29644(1) = AND(g28216, g19794)
g29969(1) = AND(g28121, g20509)
g28535(1) = AND(g11981, g27088)
g26200(2) = AND(g24688, g10678, g10658, g10627)
g25271(1) = NAND(I24462, I24463)
g26313(1) = AND(g12645, g25326)
g26082(1) = OR(g2898, g24561)
g27651(1) = AND(g22448, g25781)
g26630(1) = AND(g7592, g24419)
g27356(1) = NOR(g9429, g26657)
g28563(1) = AND(g11981, g27100)
g27369(1) = AND(g25894, g25324)
g27310(1) = AND(g26574, g23059)
I27364(1) = AND(g25541, g26424, g22698)
g27826(1) = NOR(g9501, g25821)
g27721(1) = NOR(g9672, g25805)
g27823(1) = NOR(g9792, g25805)
g30577(1) = AND(g26267, g29679)
g27765(1) = AND(g4146, g25886)
g27690(1) = AND(g25784, g23607)
g30566(1) = AND(g26247, g29507)
g28246(1) = AND(g8572, g27976)
g27299(1) = AND(g26546, g23028)
g27550(1) = NAND(g24943, g25772)
g27298(1) = AND(g26573, g23026)
g27697(1) = AND(g25785, g23649)
g27995(1) = AND(g26809, g23985)
g32040(1) = AND(g14122, g31243)
g27988(1) = AND(g26781, g23941)
g26241(2) = AND(g24688, g10678, g8778, g10627)
g27696(1) = AND(g25800, g23647)
g28547(1) = AND(g6821, g27091)
g27825(1) = NOR(g9316, g25821)
g27248(1) = OR(g24880, g25953)
g27829(1) = NOR(g7345, g25856)
g26345(1) = AND(g13051, g25505)
g26399(1) = AND(g15572, g25566)
g26652(1) = AND(g10799, g24426)
g31523(1) = AND(g7528, g29333)
g27647(1) = NOR(g3004, g26616)
g27309(1) = AND(g26603, g23057)
g27288(1) = AND(g26515, g23013)
g27659(1) = NOR(g3706, g26657)
g27379(1) = NOR(g8492, g26636)
g27343(1) = NOR(g8005, g26616)
g26541(1) = AND(g319, g24375)
g26325(1) = AND(g12644, g25370)
g26358(1) = AND(g19522, g25528)
I27349(1) = AND(g25534, g26424, g22698)
g27668(1) = AND(g1367, g25917)
g28256(1) = AND(g11398, g27984)
g27042(1) = AND(g25774, g19343)
g27771(1) = NOR(g9809, g25839)
g27678(1) = AND(g947, g25830)
g27686(1) = AND(g1291, g25849)
g26604(1) = AND(g13248, g25051)
g26395(1) = AND(g22547, g25561)
g26264(2) = AND(g24688, g8812, g8778, g10627)
g28550(1) = AND(g12009, g27092)
g27577(1) = NAND(g25019, g25002, g24988, g25765)
g26719(1) = AND(g10709, g24438)
g27879(1) = NOR(g9523, g25856)
g30670(1) = AND(g11330, g29359)
g28268(1) = AND(g8572, g27990)
g32155(1) = OR(g30935, g29475)
g27822(1) = AND(g4157, g25893)
g26389(1) = AND(g19949, g25553)
g26612(1) = AND(g901, g24407)
g26388(1) = AND(g19595, g25552)
g29381(1) = AND(g28135, g19399)
g30612(1) = AND(g26338, g29597)
g27772(1) = NOR(g7297, g25839)
g26360(1) = AND(g10589, g25533)
g26629(1) = AND(g14173, g24418)
g27344(1) = NOR(g8390, g26636)
g27733(1) = NOR(g9305, g25805)
g27665(1) = AND(g26872, g23519)
g27007(1) = NOR(g5706, g25821)
g26394(1) = AND(g22530, g25560)
g27338(1) = NOR(g9291, g26616)
g27271(1) = OR(g24547, g26053)
g27722(1) = NOR(g7247, g25805)
g31964(1) = OR(g31654, g14544)
g26190(4) = AND(g25357, g11724, g7586, g11686)
g27735(1) = NOR(g7262, g25821)
g27769(1) = NOR(g9434, g25805)
g26547(1) = AND(g13283, g25027)
g28265(1) = AND(g11367, g27989)
g31668(1) = OR(g29924, g28558)
g27664(1) = AND(g1024, g25911)
g26671(1) = AND(g316, g24429)
g27366(1) = NOR(g8016, g26636)
g31149(1) = AND(g29508, g23021)
g27931(1) = NAND(g25425, g25381, g25780)
g27674(1) = AND(g26873, g23543)
g29380(1) = AND(g28134, g19396)
g27353(1) = NOR(g8097, g26616)
g26339(1) = AND(g225, g24836)
g27704(1) = NOR(g7239, g25791)
g28236(1) = AND(g8515, g27971)
g26819(1) = AND(g106, g24490)
g27683(1) = AND(g25770, g23567)
g25215(1) = NAND(I24384, I24385)
g27244(1) = OR(g24652, g25995)
g27586(1) = NAND(g24924, g24916, g24905, g26863)
g27766(1) = NOR(g9716, g25791)
g26689(1) = AND(g15754, g24431)
g26280(1) = AND(g13051, g25248)
g27382(1) = NOR(g8219, g26657)
g26511(1) = AND(g19265, g24364)
g28537(1) = AND(g6832, g27089)
g31271(1) = AND(g29706, g23300)
g27033(1) = AND(g25767, g19273)
g26307(1) = AND(g13070, g25288)
g26670(1) = AND(g13385, g24428)
g27541(1) = AND(g26278, g23334)
g32053(1) = AND(g14176, g31509)
g31247(1) = OR(g29513, g13324)
g26487(1) = AND(g15702, g24359)
g27121(1) = AND(g136, g26326)
g31069(1) = AND(g29793, g14150)
g27682(1) = AND(g25777, g23565)
g26306(1) = AND(g13087, g25286)
g27720(1) = NOR(g9253, g25791)
g27516(1) = NOR(g9180, g26657)
g26486(1) = AND(g4423, g24358)
g27981(1) = AND(g26751, g23924)
g26223(2) = AND(g24688, g10678, g10658, g8757)
g31277(1) = OR(g29570, g28285)
g28583(1) = AND(g12009, g27112)
g26423(1) = AND(g19488, g24356)
g30936(1) = AND(g8830, g29916)
g26543(1) = AND(g12910, g24377)
g27997(1) = AND(g26813, g23995)
g26391(1) = AND(g19593, g25555)
I26948(1) = AND(g24981, g26424, g22698)
g27468(1) = NAND(g24951, g24932, g24925, g26852)
g27400(1) = NOR(g8553, g26657)
g24760(1) = NAND(I23918, I23919)
g27827(1) = NOR(g9456, g25839)
g29985(1) = AND(g28127, g20532)
g31221(1) = OR(g29494, g28204)
g26517(1) = AND(g15708, g24367)
g26362(1) = AND(g19557, g25538)
g27355(1) = NOR(g8443, g26657)
g26347(1) = AND(g262, g24850)
g29383(1) = AND(g28138, g19412)
g27367(1) = NOR(g8155, g26636)
g27345(1) = NOR(g9360, g26636)
g26351(1) = AND(g239, g24869)
g30600(1) = AND(g30287, g18975)
g27352(1) = NOR(g7975, g26616)
g26542(1) = AND(g13102, g24376)
g30607(1) = AND(g30291, g18989)
g28245(1) = AND(g11367, g27975)
g27658(1) = AND(g22491, g25786)
g31238(1) = AND(g29583, g20053)
g27732(1) = NOR(g9364, g25791)
g27878(1) = NOR(g9559, g25839)
g26381(1) = AND(g4456, g25548)
g27954(1) = NOR(g10014, g25856)
g27982(1) = NOR(g7212, g25856)
g26390(1) = AND(g4423, g25554)
g29630(1) = AND(g28212, g19781)
g30091(1) = AND(g28127, g20716)
g27479(1) = NOR(g9056, g26616)
g26397(1) = AND(g19475, g25563)
g30731(1) = AND(g11374, g29361)
g27770(1) = NOR(g9386, g25821)
g27926(1) = NOR(g9467, g25856)
g27593(1) = NAND(g24972, g24950, g24906, g26861)
g31670(1) = OR(g29937, g28573)
g26350(1) = AND(g13087, g25517)
g27027(1) = NOR(g26398, g26484)
g27287(1) = AND(g26545, g23011)
g27381(1) = NOR(g8075, g26657)
g26357(1) = AND(g22547, g25525)
g27734(1) = NOR(g9733, g25821)
g27012(1) = NOR(g6398, g25856)
g27236(1) = OR(g24620, g25974)
g24792(1) = NAND(I23950, I23951)
g26874(1) = OR(I25612, I25613)
I25908(1) = NAND(g26256, I25907)
I25909(1) = NAND(g24782, I25907)
I25244(1) = NAND(g24744, I25242)
g24380(2) = NAND(I23601, I23602)
I25221(1) = NAND(g24718, I25219)
g24369(2) = NAND(I23586, I23587)
g24802(1) = NAND(I23970, I23971)
I25220(1) = NAND(g482, I25219)
g24808(1) = NAND(I23986, I23987)
I25243(1) = NAND(g490, I25242)
I25846(1) = NAND(g26212, I25845)
I25847(1) = NAND(g24799, I25845)
g31294(1) = NOR(g11326, g29660)
g25219(1) = NOT(I24393)
g27831(1) = NOT(I26406)
g28030(1) = OR(g24018, g26874)
g31867(1) = OR(g31238, g18175)
g26881(1) = OR(g26629, g24187)
g28062(1) = OR(g27288, g21746)
g26971(1) = OR(g26325, g24333)
g26966(1) = OR(g26345, g24318)
g30390(1) = OR(g29985, g18555)
g26935(1) = NOT(I25677)
g26963(1) = OR(g26306, g24308)
g28093(1) = OR(g27981, g21951)
g26951(1) = OR(g26390, g24289)
g32978(1) = OR(g32197, g18145)
g26960(1) = OR(g26258, g24304)
g30338(1) = OR(g29613, g18240)
g26946(1) = OR(g26389, g24284)
g26891(1) = OR(g26652, g24197)
g28099(1) = OR(g27992, g22043)
g26947(1) = OR(g26394, g24285)
g30341(1) = OR(g29380, g18246)
g26892(1) = OR(g26719, g24198)
g26907(1) = OR(g26513, g24224)
g26955(1) = OR(g26391, g24293)
g26905(1) = OR(g26397, g24222)
g26901(1) = OR(g26362, g24218)
g26961(1) = OR(g26280, g24306)
g26970(1) = OR(g26308, g24332)
g26936(1) = NOT(I25680)
g31870(1) = OR(g30607, g18262)
g28098(1) = OR(g27683, g22016)
g26949(1) = OR(g26356, g24287)
g26957(1) = OR(g26517, g24295)
g26967(1) = OR(g26350, g24319)
g28102(1) = OR(g27995, g22089)
g26903(1) = OR(g26388, g24220)
g33035(1) = OR(g32019, g21872)
g28064(1) = OR(g27298, g21781)
g26959(1) = OR(g26381, g24299)
g26884(1) = OR(g26511, g24190)
g28066(1) = OR(g27553, g21819)
g26906(1) = OR(g26423, g24223)
g28068(1) = OR(g27310, g21838)
g30339(1) = OR(g29629, g18244)
g30392(1) = OR(g30091, g18558)
g26900(1) = OR(g26819, g24217)
g30347(1) = OR(g29383, g18304)
g26904(1) = OR(g26393, g24221)
g26893(1) = OR(g26753, g24199)
g26909(1) = OR(g26543, g24227)
g26890(1) = OR(g26630, g24196)
g26956(1) = OR(g26487, g24294)
g28063(1) = OR(g27541, g21773)
g26888(1) = OR(g26671, g24194)
g28105(1) = OR(g27997, g22135)
g30345(1) = OR(g29644, g18302)
g26969(1) = OR(g26313, g24329)
g31865(1) = OR(g31149, g21709)
g26883(1) = OR(g26670, g24189)
g26886(1) = OR(g26651, g24192)
g26880(1) = OR(g26610, g24186)
g26902(1) = OR(g26378, g24219)
g28095(1) = OR(g27674, g21970)
g28057(1) = OR(g27033, g18218)
g26910(1) = OR(g26571, g24228)
g26968(1) = OR(g26307, g24321)
g28082(1) = OR(g27369, g24315)
g28100(1) = OR(g27690, g22051)
g26937(1) = NOT(I25683)
g28069(1) = OR(g27564, g21865)
g31868(1) = OR(g30600, g18204)
g30391(1) = OR(g30080, g18557)
g28101(1) = OR(g27691, g22062)
g25620(1) = NOT(I24759)
g26962(1) = OR(g26295, g24307)
g26953(1) = OR(g26486, g24291)
g30340(1) = OR(g29377, g18245)
g28103(1) = OR(g27696, g22097)
g26950(1) = OR(g26357, g24288)
g25616(1) = OR(g25096, g18172)
g30389(1) = OR(g29969, g18554)
g26889(1) = OR(g26689, g24195)
g26945(1) = OR(g26379, g24283)
g30388(1) = OR(g30023, g18534)
g26911(1) = OR(g26612, g24230)
g28104(1) = OR(g27697, g22108)
g28091(1) = OR(g27665, g21913)
g28092(1) = OR(g27666, g21924)
g26948(1) = OR(g26399, g24286)
g30344(1) = OR(g29630, g18298)
g26885(1) = OR(g26541, g24191)
g28059(1) = OR(g27042, g18276)
g26908(1) = OR(g26358, g24225)
g30346(1) = OR(g29381, g18303)
g28096(1) = OR(g27988, g21997)
g26952(1) = OR(g26360, g24290)
g26954(1) = OR(g26380, g24292)
g28065(1) = OR(g27299, g21792)
g26887(1) = OR(g26542, g24193)
g25692(1) = NOT(I24839)
g26882(1) = OR(g26650, g24188)
g28097(1) = OR(g27682, g22005)
g31864(1) = OR(g31271, g21703)
g28094(1) = OR(g27673, g21959)
g28061(1) = OR(g27287, g21735)
g28067(1) = OR(g27309, g21827)
g26965(1) = OR(g26336, g24317)
g26958(1) = OR(g26395, g24297)
g26964(1) = OR(g26259, g24316)
g29385(88) = NOT(g28180)
g27700(2) = AND(g22342, g25182, g26424, g26148)
g30090(1) = NOT(g29134)
g26026(22) = NOT(I25105)
g25851(1) = NOR(g4311, g24380, g24369)
g26835(1) = NOT(I25555)
I29371(1) = NOT(g30325)
g30097(1) = NOT(g29118)
g26850(1) = NOT(I25576)
g28037(1) = NOT(g26365)
I28241(1) = NOT(g28709)
g30310(1) = NOT(g28830)
g26825(1) = NOT(I25541)
I25514(1) = NOT(g25073)
g26549(22) = NOT(I25391)
g28036(1) = NOT(g26365)
g26105(13) = NOT(I25146)
g29920(1) = NOT(g28824)
I26195(1) = NOT(g26260)
I26516(1) = NOT(g26824)
g30299(1) = NOT(g28765)
g29927(1) = NOT(g28861)
g29981(1) = NOT(g28942)
g30298(1) = OR(g28245, g27251)
g26843(1) = NOT(I25567)
g32212(3) = NOR(g8859, g31262, g11083)
g30087(1) = NOT(g29121)
g25220(1) = NOT(I24396)
g29997(1) = NOT(g29060)
g30068(1) = NOT(g29157)
g26870(1) = NOT(I25606)
g27737(1) = NOT(g26718)
g29911(1) = NOT(g28780)
g26817(1) = NOT(g25242)
g30079(1) = NOT(g29097)
g29950(1) = NOT(g28896)
g29996(1) = NOT(g28962)
g27064(8) = NOT(I25786)
g30017(1) = NOT(g29085)
g26488(22) = NOT(I25366)
g27051(5) = NOT(I25779)
g28803(8) = NOR(g27730, g22763)
g27074(8) = NOT(I25790)
g30016(1) = NOT(g29049)
g29980(1) = NOT(g28935)
I26448(1) = NOT(g26860)
g30065(1) = NOT(g29049)
I26799(1) = NOT(g27660)
g28033(1) = NOT(g26365)
I26430(1) = NOT(g26856)
g30037(1) = NOT(g29121)
I26100(1) = NOT(g26365)
g29978(1) = NOT(g28927)
g30022(1) = NOT(g29001)
g30313(1) = NOT(g28843)
g27961(1) = NOT(g26816)
g26943(1) = NOT(I25695)
g30053(1) = NOT(g29121)
g30036(1) = NOT(g29085)
g29313(1) = OR(g28284, g27270)
g25776(1) = NOR(g7166, g24380, g24369)
g27759(2) = AND(g22457, g25224, g26424, g26213)
g29923(1) = NOT(g28874)
g32137(1) = NOT(g31134)
g26941(1) = NOT(I25689)
g26519(22) = NOT(I25380)
g30074(1) = NOT(g29046)
g30931(2) = NOT(I28913)
g28032(1) = NOT(g26365)
g29942(1) = NOT(g28867)
g29993(1) = NOT(g29018)
g29965(1) = NOT(g28903)
g26576(22) = NOT(I25399)
I27238(1) = NOT(g27320)
g32192(1) = NOT(g31262)
g30052(1) = NOT(g29018)
g26400(22) = NOT(I25351)
g28120(1) = NOT(g27108)
g29922(1) = NOT(g28837)
g29953(1) = NOT(g28907)
g30100(1) = NOT(g29131)
g25771(1) = NOT(I24920)
g26862(1) = NOT(I25598)
g28126(1) = NOT(g27122)
g29983(1) = NOT(g28977)
g27724(2) = AND(g22417, g25208, g26424, g26190)
g26131(13) = NOT(I25161)
g26859(1) = NOT(I25591)
g29913(1) = NOT(g28840)
g29905(1) = NOT(g28783)
g26648(1) = NOT(g25115)
I27758(1) = NOT(g28119)
g25903(1) = NOT(I25005)
I26503(1) = NOT(g26811)
g26942(1) = NOT(I25692)
I27235(1) = NOT(g27320)
g28443(1) = NOT(I26936)
g28039(1) = NOT(g26365)
g28038(1) = NOT(g26365)
g28187(1) = NOT(I26710)
g29948(1) = NOT(g28853)
g25997(22) = NOT(I25095)
g30314(1) = OR(g28268, g27266)
g29912(1) = NOT(g28827)
I28548(1) = NOT(g28147)
g29929(1) = NOT(g28914)
I25511(1) = NOT(g25073)
g29928(1) = NOT(g28871)
g27714(2) = AND(g22384, g25195, g26424, g26171)
g30297(1) = NOT(g28758)
g29194(1) = NOT(I27492)
g27817(2) = AND(g22498, g25245, g26424, g26236)
g30088(1) = NOT(g29094)
g29999(1) = NOT(g28973)
g29998(1) = NOT(g28966)
g30311(1) = OR(g28265, g27265)
g29961(1) = NOT(g28892)
g26834(1) = NOT(I25552)
g26055(22) = NOT(I25115)
g30055(1) = NOT(g29157)
g30067(1) = NOT(g29060)
g27727(2) = AND(g22432, g25211, g26424, g26195)
g30019(1) = NOT(g29060)
g30018(1) = NOT(g28987)
g28034(1) = NOT(g26365)
g29925(1) = NOT(g28820)
g29944(1) = NOT(g28911)
g30077(1) = NOT(g29057)
g27711(2) = AND(g22369, g25193, g26424, g26166)
g30102(1) = NOT(g29157)
g27762(2) = AND(g22472, g25226, g26424, g26218)
I27677(1) = NOT(g28156)
g26510(1) = NOT(I25369)
g30076(1) = NOT(g29085)
g30085(1) = NOT(g29082)
g30054(1) = NOT(g29134)
g29995(1) = NOT(g28955)
g27414(1) = AND(g255, g26827)
g28040(1) = NOT(g26365)
g33258(1) = NOT(g32296)
g30304(1) = OR(g28255, g27259)
g28188(2) = OR(g22535, g27108)
g30039(1) = NOT(g29134)
g30306(1) = NOT(g28796)
g30038(1) = NOT(g29097)
g29960(1) = NOT(g28885)
g29955(1) = NOT(g28950)
g27832(1) = NOT(I26409)
g29967(1) = NOT(g28946)
g29994(1) = NOT(g29049)
g26851(1) = NOT(I25579)
g32138(1) = NOT(g31233)
g29977(1) = NOT(g28920)
g32424(1) = NOR(g8721, g31294)
I26508(1) = NOT(g26814)
g29976(1) = NOT(g29018)
g29893(1) = NOT(g28755)
g29939(1) = NOT(g28857)
g30063(1) = NOT(g29015)
g30021(1) = NOT(g28994)
g30300(1) = OR(g28246, g27252)
g30293(1) = OR(g28236, g27246)
g30292(1) = NOT(g28736)
g30303(1) = NOT(g28786)
g26840(1) = NOT(I25562)
g29941(1) = NOT(g28900)
g30040(1) = NOT(g29025)
g30307(1) = OR(g28256, g27260)
g33299(3) = NAND(g608, g32296, g12323)
g29906(1) = NOT(g28793)
g28194(2) = OR(g22540, g27122)
g29963(1) = NOT(g28931)
g29312(1) = NOT(g28877)
g29921(1) = NOT(g28864)
g30020(1) = NOT(g29097)
g30113(1) = NOT(g29154)
g28260(1) = AND(g27703, g26518)
g25803(1) = AND(g24798, g21024)
g28489(1) = AND(g27010, g12417)
g30003(1) = AND(g28149, g9021)
g28488(1) = AND(g27969, g17713)
g27217(1) = AND(g26236, g8418, g2610)
g29683(1) = AND(g1821, g29046)
g31962(1) = AND(g8033, g31013)
g29882(1) = AND(g2361, g29151)
g28124(1) = AND(g27368, g22842)
g29584(1) = AND(g1706, g29018)
g27186(1) = AND(g26195, g8316, g2342)
g28218(1) = AND(g27768, g26645)
g29940(1) = AND(g1740, g28758)
g29652(1) = AND(g2667, g29157)
g29804(1) = AND(g1592, g29014)
g25961(1) = AND(g25199, g20682)
g28201(1) = AND(g27499, g16720)
g28467(1) = AND(g26993, g12295)
g28494(1) = AND(g27973, g17741)
g32181(1) = AND(g31020, g19912)
g26314(8) = NOR(g24808, g24802)
g29605(1) = AND(g2445, g28973)
g32190(1) = AND(g142, g31233)
g29951(1) = AND(g1874, g28786)
g28477(1) = AND(g27966, g17676)
g29514(1) = AND(g1608, g28780)
g27493(1) = AND(g246, g26837)
g28466(1) = AND(g27960, g17637)
g32339(1) = AND(g31474, g20672)
g29535(1) = AND(g2303, g28871)
g29168(1) = OR(g27658, g26613)
g28454(1) = AND(g26976, g12233)
g32395(1) = OR(g31523, g30049)
g29649(1) = AND(g2241, g28678)
g28637(1) = AND(g22399, g27011)
g29648(1) = AND(g2112, g29121)
g29604(1) = AND(g2315, g28966)
g29563(1) = AND(g1616, g28853)
g27209(1) = AND(g26213, g8365, g2051)
g29633(1) = AND(g1978, g29085)
g29521(1) = AND(g1744, g28824)
g25989(1) = AND(g25258, g21012)
g27073(1) = AND(g7121, g3873, g3881, g26281)
g29573(1) = AND(g1752, g28892)
g29926(1) = AND(g1604, g28736)
g28139(1) = AND(g27337, g26054)
g29612(1) = AND(g27875, g28633)
g27635(9) = AND(g23032, g26281, g26424, g24996)
g28585(1) = AND(g27063, g10530)
g26994(9) = AND(g23032, g26226, g26424, g25557)
g28312(1) = AND(g27828, g26608)
g28200(1) = AND(g27652, g11383)
g29360(1) = AND(g27364, g28294)
g28115(1) = AND(g27354, g22759)
g29628(1) = AND(g27924, g28648)
g26977(9) = AND(g23032, g26261, g26424, g25550)
g28214(1) = AND(g27731, g26625)
g27040(1) = AND(g7812, g6565, g6573, g26226)
g25817(1) = AND(g24807, g21163)
g25977(1) = AND(g25236, g20875)
g32169(1) = AND(g31014, g23046)
g29645(1) = AND(g1714, g29018)
g27225(1) = OR(g2975, g26364)
g29661(1) = AND(g1687, g29015)
g29547(1) = AND(g1748, g28857)
g29895(1) = AND(g2495, g29170)
g33126(1) = AND(g9044, g32201)
g29551(1) = AND(g2173, g28867)
g29572(1) = AND(g1620, g28885)
g28273(1) = AND(g27927, g23729)
g28234(1) = AND(g27877, g26686)
g29943(1) = AND(g2165, g28765)
g29968(1) = AND(g2433, g28843)
g29855(1) = AND(g2287, g29093)
g29870(1) = AND(g2421, g29130)
g32041(1) = AND(g13913, g31262)
g29867(1) = AND(g1996, g29117)
g29894(1) = AND(g2070, g29169)
g27999(9) = AND(g23032, g26200, g26424, g25529)
g26022(1) = AND(g25271, g20751)
g32399(1) = OR(g31527, g30062)
g28240(1) = AND(g27356, g17239)
g29866(1) = AND(g1906, g29116)
g29688(1) = AND(g2509, g28713)
g29854(1) = AND(g2197, g29092)
g29511(1) = AND(g1736, g28783)
g27627(1) = AND(g13266, g25790)
g28251(1) = AND(g27826, g23662)
g28272(1) = AND(g27721, g26548)
g32034(1) = AND(g14124, g31239)
g29596(1) = AND(g27823, g28620)
g29839(1) = AND(g1728, g29045)
g29667(1) = AND(g2671, g29157)
g29838(1) = AND(g1636, g29044)
g27057(1) = AND(g7791, g6219, g6227, g26261)
g29619(1) = AND(g2269, g29060)
g32037(1) = OR(g30566, g29329)
g29601(1) = AND(g1890, g28955)
g29884(1) = AND(g2555, g29153)
g29740(1) = AND(g2648, g29154)
g29685(1) = AND(g2084, g28711)
g27161(1) = AND(g26166, g8241, g1783)
g28226(1) = AND(g27825, g26667)
g29148(1) = OR(g27651, g26606)
g28572(1) = AND(g27829, g15669)
g29964(1) = AND(g2008, g28830)
g29587(1) = AND(g2181, g28935)
g27602(9) = AND(g23032, g26244, g26424, g24966)
g29568(1) = AND(g2571, g28950)
g29638(1) = AND(g2583, g29025)
g29586(1) = AND(g1886, g28927)
g29615(1) = AND(g1844, g29049)
g28197(1) = AND(g27647, g11344)
g29684(1) = AND(g1982, g29085)
g29517(1) = AND(g1870, g28827)
g28202(1) = AND(g27659, g11413)
g29362(1) = AND(g27379, g28307)
g28111(1) = AND(g27343, g22716)
g29600(1) = AND(g1840, g29049)
g28624(1) = AND(g22357, g27009)
g28300(1) = AND(g27771, g26605)
g29530(1) = AND(g1612, g28820)
g32011(1) = AND(g8287, g31134)
g27617(9) = AND(g23032, g26264, g26424, g24982)
g28243(1) = AND(g27879, g23423)
g27467(1) = AND(g269, g26832)
g31948(1) = AND(g30670, g18884)
g29711(1) = AND(g2541, g29134)
g33252(1) = AND(g32155, g20064)
g28557(1) = AND(g27772, g15647)
g29840(1) = AND(g2153, g29056)
g29663(1) = AND(g1950, g28693)
g29553(1) = AND(g2437, g28911)
g28143(1) = AND(g27344, g26083)
g29621(1) = AND(g2449, g28994)
g29564(1) = AND(g1882, g28896)
g28217(1) = AND(g27733, g23391)
g28478(1) = AND(g27007, g12345)
g29509(1) = AND(g1600, g28755)
g29634(1) = AND(g2108, g29121)
g29851(1) = AND(g1668, g29079)
g28223(1) = AND(g27338, g17194)
g28531(1) = AND(g27722, g15608)
g33113(1) = AND(g31964, g22339)
g29574(1) = AND(g2016, g28931)
g27185(1) = AND(g26190, g8302, g1917)
g28654(1) = AND(g1030, g27108)
g29731(1) = AND(g2089, g29118)
g27439(1) = AND(g232, g26831)
g28543(1) = AND(g27735, g15628)
g28242(1) = AND(g27769, g23626)
g32094(1) = OR(g30612, g29363)
g32425(1) = AND(g31668, g21604)
g29881(1) = AND(g2040, g29150)
g28116(1) = AND(g27366, g26183)
g29662(1) = AND(g1848, g29049)
g29710(1) = AND(g2380, g29094)
I26530(1) = AND(g26365, g24096, g24097, g24098)
g28130(1) = AND(g27353, g23063)
g28523(1) = AND(g27704, g15585)
g29651(1) = AND(g2537, g29134)
g29620(1) = AND(g2399, g29097)
g25968(1) = AND(g25215, g20739)
g29646(1) = AND(g1816, g28675)
g32016(1) = AND(g8522, g31138)
g29896(1) = AND(g2599, g29171)
g32125(1) = OR(g30918, g29376)
g29582(1) = AND(g27766, g28608)
g27031(1) = OR(g26213, g26190, g26166, g26148)
g28136(1) = AND(g27382, g23135)
g29603(1) = AND(g2265, g29060)
g29549(1) = AND(g2012, g28900)
g29880(1) = AND(g1936, g29149)
g29512(1) = AND(g2161, g28793)
g32254(1) = AND(g31247, g20379)
g28673(1) = AND(g1373, g27122)
g28213(1) = AND(g27720, g23380)
g29528(1) = AND(g2429, g28874)
g28205(1) = AND(g27516, g16746)
g29869(1) = AND(g2331, g29129)
g29868(1) = AND(g2227, g29128)
g27649(1) = AND(g10820, g25820)
g29709(1) = AND(g2116, g29121)
g29708(1) = AND(g1955, g29082)
g33235(1) = OR(g32040, g30982)
g32202(1) = OR(g31069, g13410)
g32154(1) = AND(g31277, g14184)
g29602(1) = AND(g2020, g28962)
g28020(9) = AND(g23032, g26241, g26424, g25542)
g27045(1) = AND(g10295, g3171, g3179, g26244)
g29599(1) = AND(g1710, g29018)
g27032(1) = AND(g7704, g5180, g5188, g26200)
g29532(1) = AND(g1878, g28861)
g27162(1) = AND(g26171, g8259, g2208)
g29631(1) = AND(g1682, g28656)
g29364(1) = AND(g27400, g28321)
g25814(1) = AND(g24760, g13323)
g33124(1) = AND(g8945, g32296)
g28233(1) = AND(g27827, g23411)
g29687(1) = AND(g2407, g29097)
g29954(1) = AND(g2299, g28796)
g32207(1) = AND(g31221, g23323)
g27058(1) = AND(g10323, g3522, g3530, g26264)
g29525(1) = AND(g2169, g28837)
g27044(1) = AND(g7766, g5873, g5881, g26241)
g28148(1) = AND(g27355, g26093)
g29865(1) = AND(g1802, g29115)
g27146(1) = AND(g26148, g8187, g1648)
g27450(1) = OR(g2917, g26483)
g29686(1) = AND(g2246, g29057)
g28133(1) = AND(g27367, g23108)
g28229(1) = AND(g27345, g17213)
g31524(1) = AND(g29897, g20593)
g28112(1) = AND(g27352, g26162)
g29617(1) = AND(g2024, g28987)
g29984(1) = AND(g2567, g28877)
g29853(1) = AND(g1862, g29081)
g29589(1) = AND(g2575, g28977)
g29588(1) = AND(g2311, g28942)
g29524(1) = AND(g2004, g28864)
g29616(1) = AND(g1974, g29085)
g28232(1) = AND(g27732, g23586)
g28261(1) = AND(g27878, g23695)
g29642(1) = AND(g27954, g28669)
g32012(1) = AND(g8297, g31233)
g29733(1) = AND(g2675, g29157)
g28499(1) = AND(g27982, g17762)
g29665(1) = AND(g2375, g28696)
g29712(1) = AND(g2643, g28726)
g29907(1) = AND(g2629, g29177)
g28199(1) = AND(g27479, g16684)
g32173(1) = AND(g160, g31134)
g29519(1) = AND(g2295, g28840)
g31963(1) = AND(g30731, g18895)
g29637(1) = AND(g2533, g29134)
g29883(1) = AND(g2465, g29152)
g28225(1) = AND(g27770, g23400)
g28244(1) = AND(g27926, g26715)
g29577(1) = AND(g2441, g28946)
g29622(1) = AND(g2579, g29001)
g29566(1) = AND(g2307, g28907)
g31934(1) = AND(g31670, g18827)
g28010(9) = AND(g23032, g26223, g26424, g25535)
g29636(1) = AND(g2403, g29097)
g28599(1) = AND(g27027, g8922)
g29852(1) = AND(g1772, g29080)
g29664(1) = AND(g2273, g29060)
g28125(1) = AND(g27381, g26209)
g29576(1) = AND(g2177, g28903)
g29585(1) = AND(g1756, g28920)
g27037(1) = OR(g26236, g26218, g26195, g26171)
g27210(1) = AND(g26218, g8373, g2476)
g29732(1) = AND(g2514, g29131)
g28289(1) = AND(g27734, g26575)
g27039(1) = AND(g7738, g5527, g5535, g26223)
g28495(1) = AND(g27012, g12465)
g25787(1) = AND(g24792, g20887)
g29538(1) = AND(g2563, g28914)
g29496(2) = OR(g28567, g27615)
g29486(2) = OR(g28537, g27595)
g29482(2) = OR(g28524, g27588)
g27223(1) = NAND(I25908, I25909)
g27141(1) = NAND(I25846, I25847)
I26522(1) = OR(g19890, g19935, g19984, g26365)
g29495(2) = OR(g28563, g27614)
g29489(2) = OR(g28550, g27601)
g29488(2) = OR(g28547, g27600)
g29485(2) = OR(g28535, g27594)
g29501(2) = OR(g28583, g27634)
g27796(3) = NAND(g21228, g25263, g26424, g26171)
g27933(3) = NAND(g21228, g25356, g26424, g26236)
g27882(3) = NAND(g21228, g25307, g26424, g26213)
g26269(1) = NAND(I25243, I25244)
g26248(1) = NAND(I25220, I25221)
g27833(3) = NAND(g21228, g25282, g26424, g26190)
g27903(3) = NAND(g21228, g25316, g26424, g26218)
g27775(3) = NAND(g21228, g25262, g26424, g26166)
g27738(3) = NAND(g21228, g25243, g26424, g26148)
g27854(3) = NAND(g21228, g25283, g26424, g26195)
g26801(1) = NOT(I25511)
g28753(1) = NOT(I27235)
g32977(1) = OR(g32169, g21710)
g32981(1) = OR(g32425, g18206)
g33615(1) = OR(g33113, g21871)
g32979(1) = OR(g32181, g18177)
g33019(1) = OR(g32339, g18536)
g32976(1) = OR(g32207, g21704)
g32980(1) = OR(g32254, g18198)
g32985(1) = OR(g31963, g18266)
g32982(1) = OR(g31948, g18208)
g32984(1) = OR(g31934, g18264)
g31872(1) = OR(g31524, g18535)
g33538(1) = OR(g33252, g18144)
g31804(1) = NOT(g29385)
g28559(1) = NOT(g27700)
g31833(1) = NOT(g29385)
I25869(1) = NOT(g25851)
I26337(1) = NOT(g26835)
g31812(1) = NOT(g29385)
g31795(1) = NOT(I29371)
g31829(1) = NOT(g29385)
g31828(1) = NOT(g29385)
g28381(3) = NAND(g27074, g13621)
I26309(1) = NOT(g26825)
g26802(1) = NOT(I25514)
g27142(2) = NOT(g26105)
g31845(1) = NOT(g29385)
g28009(1) = NOT(I26516)
g31832(1) = NOT(g29385)
I29211(1) = NOT(g30298)
g33246(1) = NOT(g32212)
g31859(1) = NOT(g29385)
g31825(1) = NOT(g29385)
g33851(3) = NOR(g8854, g33299, g12259)
g31858(1) = NOT(g29385)
g28114(1) = AND(g25869, g27051)
g26810(1) = NOT(g25220)
g31844(1) = NOT(g29385)
I26466(1) = NOT(g26870)
I27449(1) = NOT(g27737)
g27881(1) = NOT(I26430)
g28241(1) = NOT(g27064)
g30301(1) = NOT(I28548)
g31824(1) = NOT(g29385)
I28162(1) = NOT(g28803)
I29720(1) = NOT(g30931)
g28399(1) = NOT(g27074)
I29242(1) = NOT(g29313)
I28185(1) = NOT(g28803)
g31855(1) = NOT(g29385)
g27929(1) = NOT(I26448)
g27993(1) = NOT(I26503)
g31819(1) = NOT(g29385)
g31818(1) = NOT(g29385)
g28918(1) = NOT(g27832)
g31801(1) = NOT(g29385)
g28274(4) = NOT(I26799)
I29218(1) = NOT(g30304)
I26512(1) = NOT(g26817)
I27401(1) = NOT(g27051)
g31854(1) = NOT(g29385)
I26584(1) = NOT(g26943)
I27970(1) = NOT(g28803)
I25882(1) = NOT(g25776)
g28604(1) = NOT(g27759)
I27954(1) = NOT(g28803)
g31839(1) = NOT(g29385)
g31838(1) = NOT(g29385)
g31815(1) = NOT(g29385)
I29207(1) = NOT(g30293)
I27495(1) = NOT(g27961)
g28754(1) = NOT(I27238)
I26427(1) = NOT(g26859)
g31800(1) = NOT(g29385)
g26973(2) = NOT(g26105)
g31814(1) = NOT(g29385)
I26356(1) = NOT(g26843)
g31807(1) = NOT(g29385)
I29225(1) = NOT(g30311)
g31841(1) = NOT(g29385)
g28363(3) = NAND(g27064, g13593)
g31835(1) = NOT(g29385)
I26334(1) = NOT(g26834)
I26381(1) = NOT(g26851)
g31806(1) = NOT(g29385)
I26479(1) = NOT(g25771)
I28062(1) = NOT(g29194)
I26451(1) = NOT(g26862)
g28250(1) = NOT(g27074)
g27977(2) = NOT(g26105)
g31821(1) = NOT(g29385)
I27941(1) = NOT(g28803)
g31834(1) = NOT(g29385)
g28590(1) = NOT(g27724)
g27985(2) = NOT(g26131)
g28410(3) = NAND(g27074, g13679)
g30012(2) = NOT(I28241)
g31797(1) = NOT(g29385)
g33306(3) = NAND(g776, g32212, g11679)
I27543(1) = NOT(g28187)
g29474(1) = NOT(I27758)
g28158(1) = AND(g26424, g22763, g27037)
g31796(1) = NOT(g29385)
g31840(1) = NOT(g29385)
g26990(2) = NOT(g26105)
g27155(2) = NOT(g26131)
g31847(1) = NOT(g29385)
I29717(1) = NOT(g30931)
g31851(1) = NOT(g29385)
I26581(1) = NOT(g26942)
g28406(3) = NAND(g27064, g13675)
g31820(1) = NOT(g29385)
I29228(1) = NOT(g30314)
g31846(1) = NOT(g29385)
g28395(3) = NAND(g27074, g13655)
g31827(1) = NOT(g29385)
g31803(1) = NOT(g29385)
g28391(3) = NAND(g27064, g13637)
I28174(1) = NOT(g28803)
I26130(1) = NOT(g26510)
g31826(1) = NOT(g29385)
g28579(1) = NOT(g27714)
g28615(1) = NOT(g27817)
g29317(1) = NOT(I27677)
g31811(1) = NOT(g29385)
I27927(1) = NOT(g28803)
g26987(2) = NOT(g26131)
g31850(1) = NOT(g29385)
I25743(1) = NOT(g25903)
g29186(1) = NAND(g27051, g4507)
I30904(1) = NOT(g32424)
g31802(1) = NOT(g29385)
g27698(1) = NOT(g26648)
g31857(1) = NOT(g29385)
g28376(3) = NAND(g27064, g13620)
g28593(1) = NOT(g27727)
I26578(1) = NOT(g26941)
g31856(1) = NOT(g29385)
g28575(1) = NOT(g27711)
g27004(2) = NOT(g26131)
g31831(1) = NOT(g29385)
g28606(1) = NOT(g27762)
g31843(1) = NOT(g29385)
g28326(1) = NOT(g27414)
g27972(1) = OR(g26131, g26105)
g31810(1) = NOT(g29385)
g29342(1) = NOT(g28188)
g31817(1) = NOT(g29385)
I28458(1) = NOT(g28443)
g28153(1) = AND(g26424, g22763, g27031)
g31823(1) = NOT(g29385)
I28199(1) = NOT(g28803)
g28421(3) = NAND(g27074, g13715)
I29221(1) = NOT(g30307)
g31816(1) = NOT(g29385)
g31842(1) = NOT(g29385)
g31830(1) = NOT(g29385)
g28380(1) = NOT(g27064)
g27996(1) = NOT(I26508)
g31837(1) = NOT(g29385)
g31822(1) = NOT(g29385)
g27980(1) = OR(g26105, g26131)
g31853(1) = NOT(g29385)
g31836(1) = NOT(g29385)
I29214(1) = NOT(g30300)
g31809(1) = NOT(g29385)
g31808(1) = NOT(g29385)
g27527(1) = NOT(I26195)
g31852(1) = NOT(g29385)
g27402(1) = NOT(I26100)
I26378(1) = NOT(g26850)
g31799(1) = NOT(g29385)
g31813(1) = NOT(g29385)
g33799(1) = NOT(g33299)
g29348(1) = NOT(g28194)
g31798(1) = NOT(g29385)
g31805(1) = NOT(g29385)
g31849(1) = NOT(g29385)
g31848(1) = NOT(g29385)
g31141(1) = AND(g12224, g30038)
g27410(1) = AND(g26549, g17527)
g27486(1) = AND(g26519, g17645)
g28888(1) = NAND(g27738, g8139)
g29179(1) = NOR(g9311, g28010, g7738)
g29802(1) = OR(g28243, g22871)
g27178(1) = AND(g25997, g16652)
I27529(1) = AND(g28038, g24121, g24122, g24123)
g27421(4) = AND(g8038, g26314, g9187, g9077)
g27373(1) = AND(g26488, g17477)
g28476(1) = NOR(g27627, g26547)
g27216(1) = AND(g26055, g16725)
g29107(1) = NOR(g6203, g7791, g26977)
g27117(1) = AND(g26055, g16528)
g27568(1) = AND(g26576, g17791)
g30201(1) = OR(g23412, g28557)
g33159(1) = OR(g32016, g30730)
g31788(1) = AND(g21352, g29385)
g33724(1) = AND(g14145, g33258)
g33121(1) = AND(g8748, g32212)
g28266(1) = AND(g23748, g27714)
g29183(1) = NOR(g9392, g28020, g7766)
g27416(4) = AND(g8046, g26314, g9187, g504)
g27391(1) = AND(g26549, g17505)
g27510(1) = AND(g26576, g17687)
g27489(1) = OR(g24608, g26022)
g30050(1) = AND(g22545, g28126)
g27116(1) = AND(g26026, g16527)
I27508(1) = AND(g19935, g24082, g24083, g28033)
g27395(4) = AND(g8046, g26314, g9187, g9077)
g27430(1) = AND(g26488, g17579)
g27517(1) = AND(g26400, g17707)
g29344(1) = AND(g29168, g18932)
g28481(1) = NOR(g3506, g10323, g27617)
g27130(1) = AND(g26026, g16585)
g29144(1) = NOR(g9518, g26977)
g27523(1) = AND(g26549, g17718)
g27222(1) = AND(g26055, g13932)
g27494(4) = AND(g8038, g26314, g518, g9077)
g27437(1) = AND(g26576, g17589)
g27135(1) = OR(g24387, g25803)
g27347(1) = AND(g26400, g17390)
g33099(1) = AND(g32395, g18944)
g31777(1) = AND(g21343, g29385)
g27372(1) = AND(g26488, g17476)
g27137(1) = AND(g26026, g16606)
g31140(1) = AND(g2102, g30037)
g29165(1) = NOR(g5881, g28020)
g27273(1) = NAND(g10504, g26131, g26105)
g29007(1) = NOR(g9269, g28010)
g29071(1) = NOR(g5873, g28020)
g27436(1) = AND(g26576, g17588)
g27346(1) = AND(g26400, g17389)
g31776(1) = AND(g21329, g29385)
g31147(1) = AND(g12286, g30054)
g27153(1) = AND(g26055, g16629)
g28965(1) = NAND(g27882, g8255)
g27409(1) = AND(g26519, g17524)
g27136(1) = AND(g26026, g16605)
g27408(1) = AND(g26519, g17523)
g31151(1) = AND(g10037, g30065)
g29106(1) = NOR(g9451, g28020)
g29175(1) = NOR(g6227, g26977)
g27474(4) = AND(g8038, g26314, g518, g504)
g27537(1) = AND(g26549, g17742)
g29904(1) = OR(g28312, g26146)
I27513(1) = AND(g19984, g24089, g24090, g28034)
g27445(4) = AND(g8038, g26314, g9187, g504)
g31472(1) = OR(g29642, g28352)
g31120(1) = AND(g1700, g29976)
g31146(1) = AND(g12285, g30053)
g29035(1) = NOR(g9321, g28020)
g28552(1) = NOR(g10295, g27602)
g29734(1) = OR(g28201, g15872)
g27390(1) = AND(g26549, g17504)
g27522(1) = AND(g26549, g17717)
g27483(1) = AND(g26488, g17642)
g29768(1) = OR(g22760, g28229)
g27536(1) = AND(g26519, g17738)
g29786(1) = OR(g22843, g28240)
g30176(1) = OR(g23392, g28531)
g27183(1) = AND(g26055, g16658)
g27469(4) = AND(g8046, g26314, g518, g9077)
g27508(1) = AND(g26549, g17684)
g27213(1) = AND(g26026, g16721)
g29879(1) = OR(g28289, g26096)
g27452(1) = AND(g26400, g17600)
g28899(1) = NAND(g27833, g14612)
g31211(1) = AND(g10156, g30102)
g27282(1) = NAND(g11192, g26269, g26248, g479)
g31375(1) = OR(g29628, g28339)
g28263(1) = AND(g23747, g27711)
g27413(1) = AND(g26576, g17530)
g29142(1) = NOR(g5535, g28010)
g29198(1) = NOR(g7766, g28020)
g27113(1) = AND(g25997, g16522)
g30081(1) = OR(g28454, g11366)
g27357(1) = AND(g26400, g17414)
g27105(1) = AND(g26026, g16511)
g29484(1) = OR(g28124, g22191)
g28514(1) = NOR(g8165, g27617)
g31150(1) = AND(g1682, g30063)
g29481(1) = OR(g28117, g28125)
g29145(1) = NOR(g6549, g7812, g26994)
g29480(1) = OR(g28115, g22172)
g27482(1) = AND(g26488, g17641)
g28945(1) = NAND(g27854, g8211)
g27440(4) = AND(g8046, g26314, g518, g504)
g27204(1) = AND(g26026, g16689)
g28462(1) = NOR(g3512, g27617)
g29717(1) = OR(g28200, g10883)
g27090(1) = AND(g25997, g16423)
g33102(1) = AND(g32399, g18978)
g29483(1) = OR(g25801, g28130)
g28468(1) = NOR(g3155, g10295, g27602)
g27505(1) = AND(g26519, g17681)
g27404(1) = AND(g26400, g17518)
g30127(1) = OR(g28494, g16805)
g27212(1) = AND(g25997, g16717)
g28938(1) = NAND(g27796, g8205)
g27149(1) = AND(g25997, g16623)
g27433(1) = AND(g26519, g17583)
g27387(1) = AND(g26488, g17499)
g27148(1) = AND(g25997, g16622)
g27104(1) = AND(g25997, g16510)
g29034(1) = NOR(g5527, g28010)
g29191(1) = NOR(g7738, g28010)
g28491(1) = NOR(g8114, g27617)
g27412(1) = AND(g26576, g17529)
g27229(1) = AND(g26055, g16774)
g27228(1) = AND(g26055, g16773)
g31131(1) = AND(g2393, g30020)
g31210(1) = AND(g2509, g30100)
g29716(1) = OR(g28199, g15856)
g27386(1) = AND(g26488, g17498)
g27096(1) = AND(g26026, g16475)
g28990(1) = NAND(g27882, g8310)
g29005(1) = NOR(g5164, g7704, g27999)
g31187(1) = AND(g10118, g30090)
g27428(1) = AND(g26400, g17576)
g29506(1) = OR(g28148, g25880)
g27549(1) = AND(g26576, g14785)
g31169(1) = AND(g10083, g30079)
g27548(1) = AND(g26576, g17763)
g31168(1) = AND(g2241, g30077)
g27504(1) = AND(g26519, g17680)
g29764(1) = OR(g28219, g28226)
g29476(1) = OR(g28108, g28112)
g29777(1) = OR(g28227, g28234)
g31319(1) = OR(g29612, g28324)
g27129(1) = AND(g26026, g16584)
g27128(1) = AND(g25997, g16583)
g28870(1) = NAND(g27796, g14588)
g31186(1) = AND(g2375, g30088)
g33186(1) = AND(g32037, g22830)
g28986(1) = NOR(g5517, g28010)
g28980(1) = NAND(g27933, g14680)
g27432(1) = AND(g26519, g17582)
g28519(1) = NOR(g8011, g27602, g10295)
g27461(1) = AND(g26576, g17611)
g31123(1) = AND(g1834, g29994)
g28290(1) = AND(g23780, g27759)
g27650(1) = AND(g26519, g15479)
g29033(1) = NOR(g5511, g7738, g28010)
g27132(1) = AND(g26055, g16589)
g29334(1) = AND(g29148, g18908)
I27524(1) = AND(g28037, g24114, g24115, g24116)
g30093(1) = OR(g28467, g11397)
g27375(1) = AND(g26519, g17479)
g29791(1) = OR(g28233, g22859)
g29028(1) = NAND(g27933, g8381)
g31142(1) = AND(g2527, g30039)
g29849(1) = OR(g26049, g28273)
g29173(1) = NOR(g9259, g27999, g7704)
g27459(1) = AND(g26549, g17609)
g28510(1) = NOR(g3530, g27617)
g29181(1) = NOR(g6573, g26994)
g31130(1) = AND(g12191, g30019)
g27545(1) = AND(g26519, g17756)
g29012(1) = NOR(g5863, g28020)
g28856(1) = NAND(g27738, g8093)
g29756(1) = OR(g22717, g28223)
g28457(1) = NOR(g7980, g27602)
g31222(1) = AND(g2643, g30113)
g29193(1) = NOR(g9529, g26994, g7812)
g28521(1) = NOR(g27649, g26604)
g31790(1) = AND(g21299, g29385)
g29848(1) = OR(g28260, g26077)
g33291(1) = OR(g32154, g13477)
I27519(1) = AND(g28036, g24107, g24108, g24109)
g31209(1) = AND(g2084, g30097)
g29189(1) = NOR(g9462, g26977, g7791)
g28930(1) = NAND(g27833, g8201)
g27374(1) = AND(g26519, g17478)
g31122(1) = AND(g12144, g29993)
g33122(1) = AND(g8859, g32192)
g27669(1) = AND(g26840, g13278)
g29735(1) = OR(g28202, g10898)
g31153(1) = AND(g12336, g30068)
g27392(1) = AND(g26576, g17507)
g27559(1) = AND(g26576, g17777)
g27525(1) = AND(g26576, g17720)
g27488(1) = AND(g26549, g17648)
g27558(1) = AND(g26576, g17776)
g28895(1) = NAND(g27775, g8146)
g28280(1) = AND(g23761, g27724)
I27539(1) = AND(g28040, g24135, g24136, g24137)
g27460(1) = AND(g26549, g17610)
g29790(1) = OR(g25975, g28242)
g29164(1) = NOR(g9444, g28010)
g27267(1) = AND(g26026, g17124)
g28860(1) = NAND(g27775, g14586)
g29069(1) = NOR(g9381, g28010)
g30103(1) = OR(g28477, g16731)
g28509(1) = NOR(g8107, g27602)
g28470(1) = NOR(g8021, g27617)
g27219(1) = AND(g26026, g16742)
g27218(1) = AND(g25997, g16740)
g28520(1) = NOR(g8229, g27635)
g27455(1) = AND(g26488, g17603)
g28910(1) = NAND(g27854, g14614)
g27201(1) = AND(g25997, g16685)
g29070(1) = NOR(g5857, g7766, g28020)
g28976(1) = NAND(g27903, g8273)
g28480(1) = NOR(g8059, g27602)
g29200(1) = NOR(g7791, g26977)
g29813(1) = OR(g26020, g28261)
g27118(1) = AND(g26055, g16529)
g29072(1) = NOR(g9402, g26977)
g28923(1) = NAND(g27775, g8195)
g30061(1) = AND(g1036, g28188)
g27177(1) = AND(g25997, g16651)
g30114(1) = OR(g28488, g16761)
g30163(1) = OR(g23381, g28523)
g28969(1) = NAND(g27854, g8267)
g31152(1) = AND(g10039, g30067)
g29184(1) = NOR(g9631, g26994)
g27485(1) = AND(g26519, g17644)
g27431(1) = OR(g24582, g25977)
g31307(1) = OR(g29596, g28311)
g27454(1) = AND(g26488, g17602)
g31787(1) = AND(g21281, g29385)
g27519(1) = AND(g26488, g17710)
g33105(1) = AND(g26298, g32138)
g27518(1) = AND(g26488, g17709)
g27154(1) = AND(g26055, g16630)
g30141(1) = OR(g28499, g16844)
g28469(1) = NOR(g3171, g27602)
g28106(1) = NOR(g7812, g26994)
g28492(1) = NOR(g3857, g7121, g27635)
g29180(1) = NOR(g9569, g26977)
g29174(1) = NOR(g9511, g28020)
g27215(1) = AND(g26055, g16724)
g27501(1) = AND(g26400, g17673)
g27348(1) = AND(g26488, g17392)
g31778(1) = AND(g21369, g29385)
g30189(1) = OR(g23401, g28543)
g27139(1) = AND(g26055, g16608)
g27653(1) = AND(g26549, g15562)
g27138(1) = AND(g26055, g16607)
g33233(1) = AND(g32094, g23005)
g28498(1) = NOR(g8172, g27635)
g28414(1) = NOR(g27467, g26347)
g27115(1) = AND(g26026, g16526)
g33723(1) = AND(g14091, g33299)
g28035(1) = AND(g24103, I26530, I26531)
g31148(1) = AND(g2661, g30055)
g33104(1) = AND(g26296, g32137)
g28934(1) = NAND(g27882, g14641)
g27214(1) = AND(g26026, g13901)
g27207(1) = AND(g26055, g16692)
g27539(1) = AND(g26576, g17745)
g31293(1) = OR(g29582, g28299)
g27538(1) = AND(g26549, g14744)
g29146(1) = NOR(g6565, g26994)
g28253(1) = AND(g23719, g27700)
g27407(1) = AND(g26488, g17522)
I27534(1) = AND(g28039, g24128, g24129, g24130)
g30128(1) = OR(g28495, g11497)
g28209(1) = OR(g27223, g27141)
g29167(1) = NOR(g9576, g26994)
g27405(1) = OR(g24572, g25968)
g29370(1) = NOR(g28585, g28599)
g27582(1) = NAND(g10857, g26131, g26105)
g27206(1) = AND(g26055, g16691)
g28340(1) = NOR(g27439, g26339)
g27114(1) = AND(g25997, g16523)
g31129(1) = AND(g1968, g30017)
g27435(1) = AND(g26549, g17585)
g27107(1) = AND(g26055, g16514)
g27383(1) = OR(g24569, g25961)
g31128(1) = AND(g12187, g30016)
g33245(1) = AND(g32125, g19961)
g28493(1) = NOR(g3873, g27635)
g28292(1) = AND(g23781, g27762)
g28953(1) = NOR(g5170, g27999)
g27406(1) = AND(g26488, g17521)
g27361(1) = AND(g26519, g17419)
g31001(1) = OR(g29360, g28151)
g27500(1) = AND(g26400, g17672)
g27221(1) = AND(g26055, g16747)
g33794(1) = OR(g33126, g32053)
g29801(1) = OR(g25987, g28251)
g27106(1) = AND(g26026, g16512)
g27371(1) = AND(g26400, g17473)
g27234(1) = AND(g26055, g16814)
g28584(1) = NOR(g7121, g27635)
g31145(1) = AND(g9970, g30052)
g28958(1) = NAND(g27833, g8249)
g27507(1) = AND(g26549, g17683)
g30279(1) = OR(g28637, g27668)
g29504(1) = OR(g28143, g25875)
g27359(1) = AND(g26488, g17416)
g29754(1) = OR(g28215, g28218)
g27535(1) = AND(g26519, g17737)
g27434(1) = AND(g26549, g17584)
g27358(1) = AND(g26400, g17415)
g27159(1) = OR(g25814, g12953)
g33244(1) = AND(g32190, g23152)
g29006(1) = NOR(g5180, g27999)
g28540(1) = NOR(g8125, g27635, g7121)
g29187(1) = NOR(g7704, g27999)
g27134(1) = AND(g25997, g16602)
g30214(1) = OR(g23424, g28572)
g31007(1) = OR(g29364, g28159)
g28949(1) = NAND(g27903, g14643)
g27491(1) = AND(g26576, g17652)
g33817(1) = AND(g33235, g20102)
g33322(1) = AND(g32202, g20450)
g29502(1) = OR(g28139, g25871)
g29040(1) = NOR(g6209, g26977)
g27262(1) = AND(g25997, g17092)
g27521(1) = AND(g26519, g14700)
g29479(1) = OR(g28113, g28116)
g27389(1) = AND(g26519, g17503)
g27388(1) = AND(g26519, g17502)
g28282(1) = AND(g23762, g27727)
g27534(1) = AND(g26488, g17735)
g28302(1) = AND(g23809, g27817)
g27272(1) = AND(g26055, g17144)
I27503(1) = AND(g19890, g24075, g24076, g28032)
g27462(1) = AND(g26576, g17612)
g28823(1) = NAND(g27738, g14565)
g30104(1) = OR(g28478, g11427)
g29748(1) = OR(g28210, g28214)
g28515(1) = NOR(g3881, g27635)
g27360(1) = AND(g26488, g17417)
g29892(1) = OR(g28300, g26120)
g29478(1) = OR(g28111, g22160)
g27152(1) = OR(g24393, g25817)
g27451(1) = AND(g26400, g17599)
g27220(1) = AND(g26026, g16743)
g27628(1) = AND(g26400, g18061)
g28452(1) = NOR(g3161, g27602)
g29692(1) = OR(g28197, g10873)
g27370(1) = AND(g26400, g17472)
g31124(1) = AND(g2259, g29997)
g27151(1) = AND(g26026, g16626)
g29141(1) = NOR(g9374, g27999)
g27227(1) = AND(g26026, g16771)
g27540(1) = AND(g26576, g17746)
g30035(1) = AND(g22539, g28120)
g27203(1) = AND(g26026, g16688)
g29753(1) = OR(g28213, g22720)
g29792(1) = OR(g28235, g28244)
g27645(1) = AND(g26488, g15344)
g28483(1) = NOR(g8080, g27635)
g29032(1) = NOR(g9300, g27999)
g27427(1) = AND(g26400, g17575)
g27126(1) = OR(g24378, g25787)
g27661(1) = AND(g26576, g15568)
g27547(1) = AND(g26549, g17759)
g31167(1) = AND(g10080, g30076)
g27481(1) = AND(g26400, g14630)
g29763(1) = OR(g28217, g22762)
g29490(1) = OR(g25832, g28136)
g27127(1) = AND(g25997, g16582)
g27490(1) = AND(g26576, g17651)
g27376(1) = AND(g26549, g17481)
g27385(1) = AND(g26400, g17497)
g29741(1) = OR(g28205, g15883)
g27103(1) = AND(g25997, g16509)
g27095(1) = AND(g25997, g16473)
g27181(1) = AND(g26026, g16655)
g28475(1) = NOR(g3863, g27635)
g28496(1) = NOR(g3179, g27602)
g27520(1) = AND(g26519, g17714)
g30073(1) = AND(g1379, g28194)
g27546(1) = AND(g26549, g17758)
g31166(1) = AND(g1816, g30074)
g27211(1) = AND(g25997, g16716)
g29776(1) = OR(g28225, g22846)
g29077(1) = NOR(g6555, g26994)
g28425(1) = NOR(g27493, g26351)
g27339(1) = AND(g26400, g17308)
g29864(1) = OR(g28272, g26086)
g31185(1) = AND(g10114, g30087)
g27411(1) = AND(g26549, g17528)
g27503(1) = AND(g26488, g14668)
g27202(1) = AND(g25997, g13876)
g29004(1) = NAND(g27933, g8330)
g27384(1) = AND(g26400, g17496)
g27094(1) = AND(g25997, g16472)
g28529(1) = NOR(g8070, g27617, g10323)
g31139(1) = AND(g12221, g30036)
g27526(1) = AND(g26576, g17721)
g28906(1) = NAND(g27796, g8150)
g27457(1) = AND(g26519, g17606)
g30564(1) = AND(g21358, g29385)
g29775(1) = OR(g25966, g28232)
g29487(1) = OR(g25815, g28133)
g31184(1) = AND(g1950, g30085)
g33232(1) = OR(g32034, g30936)
g29109(1) = NOR(g9472, g26994)
g30270(1) = OR(g28624, g27664)
g27480(1) = AND(g26400, g17638)
g28997(1) = NAND(g27903, g8324)
g33241(1) = AND(g32173, g23128)
g28482(1) = NOR(g3522, g27617)
g28568(1) = NOR(g10323, g27617)
g27180(1) = AND(g26026, g16654)
g27131(1) = AND(g26055, g16588)
g29108(1) = NOR(g6219, g26977)
g28981(1) = NOR(g9234, g27999)
g31002(1) = OR(g29362, g28154)
g27502(1) = AND(g26488, g17677)
g27557(1) = AND(g26549, g17774)
g27458(1) = OR(g24590, g25989)
g31759(1) = AND(g21291, g29385)
g33123(1) = OR(g31962, g30577)
g30115(1) = OR(g28489, g11449)
g30092(1) = OR(g28466, g16699)
g29104(1) = NOR(g5188, g27999)
I26643(1) = OR(g27073, g27058, g27045, g27040)
g28191(1) = OR(g27217, g27210, g27186, g27162)
I26644(1) = OR(g27057, g27044, g27039, g27032)
g28186(1) = OR(g27209, g27185, g27161, g27146)
g28031(1) = NOR(g21209, I26522, I26523)
I26459(2) = NAND(g26576, g14306)
I29295(2) = NAND(g29495, g12117)
I26093(2) = NAND(g26055, g13539)
I26417(2) = NAND(g26519, g14247)
I29313(2) = NAND(g29501, g12154)
g28109(1) = NAND(g27051, g25783)
I26438(2) = NAND(g26549, g14271)
I29269(2) = NAND(g29486, g12050)
I29277(2) = NAND(g29488, g12081)
I29284(2) = NAND(g29489, g12085)
I26049(2) = NAND(g25997, g13500)
g28131(1) = NAND(g27051, g25838)
I29253(2) = NAND(g29482, g12017)
I26393(2) = NAND(g26488, g14227)
I29302(2) = NAND(g29496, g12121)
I26070(2) = NAND(g26026, g13517)
I26366(2) = NAND(g26400, g14211)
I29261(2) = NAND(g29485, g12046)
g32185(1) = NOT(I29717)
g32454(1) = OR(g30322, g31795)
g33535(1) = OR(g33233, g21711)
g33539(1) = OR(g33245, g18178)
g33537(1) = OR(g33244, g21716)
g33534(1) = OR(g33186, g21700)
g30337(1) = OR(g29334, g18220)
g28080(1) = NOT(I26581)
g28079(1) = NOT(I26578)
g30343(1) = OR(g29344, g18278)
g33536(1) = OR(g33241, g21715)
g29209(1) = NOT(I27543)
g33540(1) = OR(g33099, g18207)
g33964(1) = OR(g33817, g18146)
g33608(1) = OR(g33322, g18537)
g33542(1) = OR(g33102, g18265)
g28081(1) = NOT(I26584)
g29722(2) = NAND(g28410, g13742)
g29719(2) = NAND(g28406, g13739)
g30217(1) = NOT(I28458)
g29812(1) = NOT(g28381)
g27880(1) = NOT(I26427)
I29182(1) = NOT(g30012)
g27967(1) = NOT(I26479)
g27773(1) = NOT(I26378)
I28002(1) = NOT(g28153)
g29672(2) = NAND(g28376, g13672)
g34161(1) = NOT(g33851)
I28434(1) = NOT(g28114)
g27930(1) = NOT(I26451)
g29147(1) = NOT(I27449)
I27368(1) = NOT(g27881)
g29029(2) = AND(g14506, g25227, g26424, g27494)
I28832(1) = NOT(g30301)
g28959(2) = AND(g17401, g25194, g26424, g27440)
g32186(1) = NOT(I29720)
g31658(6) = NOT(I29242)
g29956(2) = NOT(I28185)
g27708(1) = NOT(I26334)
I27232(1) = NOT(g27993)
g27928(1) = NOT(g26810)
I26952(1) = NOT(g27972)
g30218(1) = NOT(g28918)
g29339(2) = NOT(g28274)
g27998(1) = NOT(I26512)
g31624(6) = NOT(I29218)
I28572(1) = NOT(g28274)
g29067(1) = NOT(I27401)
g28939(2) = AND(g17321, g25184, g26424, g27421)
g29689(2) = NOT(I27954)
g30142(1) = NOT(g28754)
g29930(2) = NOT(I28162)
g31601(6) = NOT(I29207)
g27774(1) = NOT(I26381)
I26880(1) = NOT(g27527)
g28970(2) = AND(g17405, g25196, g26424, g27445)
g27675(1) = NOT(I26309)
g29737(2) = NAND(g28421, g13779)
g28652(1) = AND(g27282, g10288)
g27736(1) = NOT(I26356)
g31639(6) = NOT(I29225)
g29800(1) = NOT(g28363)
g27709(1) = NOT(I26337)
g29814(19) = NOT(I28062)
g27013(1) = NOT(I25743)
g29863(1) = NOT(g28410)
g33797(1) = NOT(g33306)
g27830(1) = NOT(g26802)
I27314(1) = NOT(g28009)
I28579(1) = NOT(g29474)
I28014(1) = NOT(g28158)
g29505(1) = NOT(g29186)
I29185(1) = NOT(g30012)
g27956(1) = NOT(I26466)
g29676(2) = NAND(g28381, g13676)
g29702(2) = NAND(g28395, g13712)
g29862(1) = NOT(g28406)
g29847(1) = NOT(g28395)
I28851(1) = NOT(g29317)
g33823(3) = NOR(g8774, g33306, g11083)
g29694(2) = NAND(g28391, g13709)
g28998(2) = AND(g17424, g25212, g26424, g27474)
g30318(2) = NOT(g28274)
g29846(1) = NOT(g28391)
g29675(1) = NOR(g28380, g8236, g8354)
g27438(1) = NOT(I26130)
g29945(2) = NOT(I28174)
g31646(6) = NOT(I29228)
g28889(2) = AND(g17292, g25169, g26424, g27395)
g30286(1) = OR(g28191, g28186)
g33378(1) = NOT(I30904)
I27388(1) = NOT(g27698)
g29811(1) = NOT(g28376)
I26929(1) = NOT(g27980)
g28991(2) = AND(g14438, g25209, g26424, g27469)
g27163(13) = NOT(I25869)
g28140(1) = OR(I26643, I26644)
I27391(1) = NOT(g27929)
g29970(2) = NOT(I28199)
g29878(1) = NOT(g28421)
g31631(6) = NOT(I29221)
I27253(1) = NOT(g27996)
g29669(2) = NOT(I27941)
g29195(1) = NOT(I27495)
g29657(2) = NAND(g28363, g13634)
g29713(2) = NOT(I27970)
g34174(3) = NAND(g617, g33851, g12323)
g31616(6) = NOT(I29214)
g29705(1) = NOR(g28399, g8284, g8404)
g31609(6) = NOT(I29211)
g29653(2) = NOT(I27927)
g28924(2) = AND(g17317, g25183, g26424, g27416)
g27187(13) = NOT(I25882)
g28743(1) = OR(g27517, g16758)
g28322(1) = OR(g27117, g15809)
g28670(1) = OR(g27412, g16618)
g32217(1) = OR(g31129, g29616)
g32257(1) = OR(g31184, g29708)
g29515(1) = AND(g28888, g22342)
g29991(1) = AND(g29179, g12922)
g31500(1) = AND(g29802, g23449)
g28720(1) = OR(g27486, g16704)
g29206(1) = AND(g24124, I27528, I27529)
g28308(1) = OR(g27105, g15795)
g28267(1) = AND(g7328, g2227, g27421)
g28306(1) = OR(g27104, g15794)
g30026(1) = AND(g28476, g25064)
g28687(1) = OR(g27434, g16638)
g29345(1) = AND(g4749, g28376)
g29332(1) = AND(g29107, g22170)
g31541(1) = AND(g22536, g29348)
g31789(1) = AND(g30201, g24013)
g33789(1) = AND(g33159, g23022)
g32249(1) = OR(g31169, g29687)
g28716(1) = OR(g27481, g13887)
g32228(1) = OR(g31147, g29651)
g28715(1) = OR(g27480, g16700)
g30011(1) = AND(g29183, g12930)
g28588(1) = AND(g27489, g20499)
g28344(1) = OR(g27136, g15820)
g28254(1) = AND(g7268, g1668, g27395)
g28270(1) = NAND(g10504, g26105, g26987)
g28335(1) = OR(g27132, g15818)
g30002(1) = AND(g28481, g23487)
g30057(1) = AND(g29144, g9462)
g31772(1) = OR(g30035, g28654)
g28733(1) = OR(g27507, g16735)
g28309(1) = OR(g27106, g15796)
g28719(1) = OR(g27485, g16703)
g28239(1) = AND(g27135, g19659)
g28772(1) = OR(g27534, g16802)
g28320(1) = OR(g27116, g15808)
g30056(1) = AND(g29165, g12659)
g28317(1) = OR(g27114, g15805)
g28342(1) = OR(g27134, g15819)
g28375(1) = OR(g27183, g15851)
g28439(1) = AND(g27273, g10233)
g28428(1) = OR(g27227, g15912)
g29990(1) = AND(g29007, g9239)
g30031(1) = AND(g29071, g10540)
g28664(1) = OR(g27408, g16613)
g28512(1) = NAND(g10857, g27155, g27142)
g28662(1) = OR(g27407, g16612)
g28390(1) = OR(g27207, g15861)
g32243(1) = OR(g31166, g29683)
g29534(1) = AND(g28965, g22457)
g28705(1) = OR(g27460, g16672)
g31779(1) = OR(g30050, g28673)
g28751(1) = OR(g27526, g16766)
g32271(1) = OR(g31209, g29731)
g30043(1) = AND(g29106, g9392)
g28732(1) = OR(g27505, g16734)
g30069(1) = AND(g29175, g12708)
g28316(1) = OR(g27113, g15804)
g28400(1) = OR(g27211, g15870)
g31540(1) = AND(g29904, g23548)
g28799(3) = AND(g21434, g26424, g25348, g27445)
g32341(1) = AND(g31472, g23610)
g30010(1) = AND(g29035, g9274)
g29591(1) = AND(g28552, g11346)
g28332(1) = OR(g27130, g15815)
g31290(1) = AND(g29734, g23335)
g28761(3) = AND(g21434, g26424, g25299, g27416)
g28388(1) = OR(g27204, g15859)
g28387(1) = OR(g27203, g15858)
g28374(1) = OR(g27181, g15850)
g31481(1) = AND(g29768, g23417)
g31490(1) = AND(g29786, g23429)
g29203(1) = AND(g24095, I27513, I27514)
g31784(1) = AND(g30176, g24003)
g28430(1) = OR(g27229, g15914)
g28884(1) = OR(g27568, g16885)
g28704(1) = OR(g27459, g16671)
g31520(1) = AND(g29879, g23507)
g29632(1) = AND(g28899, g22417)
g32221(1) = OR(g31140, g29634)
g32334(1) = AND(g31375, g23568)
g32220(1) = OR(g31139, g29633)
g28331(1) = OR(g27129, g15814)
g29354(1) = AND(g4961, g28421)
g28418(1) = OR(g27220, g15882)
g30042(1) = AND(g29142, g12601)
g28748(1) = OR(g27522, g16763)
g28833(3) = AND(g21434, g26424, g25388, g27469)
g28644(1) = OR(g27387, g16593)
g30030(1) = AND(g29198, g12347)
g28776(1) = OR(g27538, g13974)
g31707(1) = AND(g30081, g23886)
g28698(1) = OR(g27451, g16666)
g28389(1) = OR(g27206, g15860)
g31067(1) = AND(g29484, g22868)
g29625(1) = AND(g28514, g14226)
g31019(1) = AND(g29481, g22856)
g29338(1) = AND(g29145, g22181)
g28817(1) = OR(g27548, g16845)
g31018(1) = AND(g29480, g22855)
g31526(1) = AND(g22521, g29342)
g29527(1) = AND(g28945, g22432)
g28789(3) = AND(g21434, g26424, g25340, g27440)
g28775(1) = OR(g27537, g16806)
g29581(1) = AND(g28462, g11796)
g31280(1) = AND(g29717, g23305)
g28622(1) = OR(g27360, g16519)
g28651(1) = OR(g27392, g16599)
g29202(1) = AND(g24088, I27508, I27509)
g28291(1) = AND(g7411, g2070, g27469)
g29590(1) = AND(g2625, g28615)
g31066(1) = AND(g29483, g22865)
g29986(1) = AND(g28468, g23473)
g28179(1) = OR(g27494, g27474, g27445, g27421)
g31763(1) = AND(g30127, g23965)
g28405(1) = OR(g27216, g15875)
g28747(1) = OR(g27521, g13942)
g28631(1) = OR(g27372, g16534)
g29526(1) = AND(g28938, g22384)
g28621(1) = OR(g27359, g16518)
g30009(1) = AND(g29034, g10518)
g30008(1) = AND(g29191, g12297)
g32223(1) = OR(g31142, g29637)
g29624(1) = AND(g28491, g8070)
g28728(1) = OR(g27501, g16730)
g28404(1) = OR(g27215, g15874)
g28416(1) = OR(g27218, g15880)
g28727(1) = OR(g27500, g16729)
g28640(1) = OR(g27384, g16590)
g28611(1) = OR(g27348, g16485)
g31278(1) = AND(g29716, g23302)
g29550(1) = AND(g28990, g22457)
g29314(1) = AND(g29005, g22144)
g28690(1) = OR(g27436, g16641)
g31143(1) = AND(g29506, g22999)
g28203(1) = NAND(g12546, g27985, g27977)
g28852(1) = OR(g27559, g16871)
g34125(1) = OR(g33724, g33124)
g32262(1) = OR(g31186, g29710)
g31478(1) = AND(g29764, g23410)
g31015(1) = AND(g29476, g22758)
g31486(1) = AND(g29777, g23422)
g32327(1) = AND(g31319, g23544)
g29618(1) = AND(g28870, g22384)
g29975(1) = AND(g28986, g10420)
g28665(1) = OR(g27409, g16614)
g32219(1) = OR(g31131, g29620)
g29666(1) = AND(g28980, g22498)
g28281(1) = AND(g7362, g1936, g27440)
g28739(3) = AND(g21434, g26424, g25274, g27395)
g29580(1) = AND(g28519, g14186)
g29321(1) = AND(g29033, g22148)
g29531(1) = AND(g1664, g28559)
g28680(1) = OR(g27427, g16633)
g28230(1) = OR(g27669, g14261)
g28729(1) = OR(g27502, g16732)
g28298(1) = NAND(g10533, g26131, g26990)
g28723(1) = OR(g27490, g16706)
g28435(1) = OR(g27234, g15967)
g31746(1) = AND(g30093, g23905)
g31493(1) = AND(g29791, g23434)
g29569(1) = AND(g29028, g22498)
g28286(1) = OR(g27090, g15757)
g32222(1) = OR(g31141, g29636)
g31517(1) = AND(g29849, g23482)
g28297(1) = OR(g27096, g15785)
g28359(1) = OR(g27151, g15838)
g28323(1) = OR(g27118, g15810)
g29974(1) = AND(g29173, g12914)
g29639(1) = AND(g28510, g11618)
g30082(1) = AND(g29181, g12752)
g32259(1) = OR(g31185, g29709)
g28371(1) = OR(g27177, g15847)
g29992(1) = AND(g29012, g10490)
g29510(1) = AND(g28856, g22342)
g31475(1) = AND(g29756, g23406)
g29579(1) = AND(g28457, g7964)
g29578(1) = AND(g2491, g28606)
g29835(1) = AND(g28326, g24866)
g28773(1) = OR(g27535, g16803)
g32236(1) = OR(g31152, g29664)
g32285(1) = OR(g31222, g29740)
g30048(1) = AND(g29193, g12945)
g30004(1) = AND(g28521, g25837)
g28700(1) = OR(g27454, g16668)
g31516(1) = AND(g29848, g23476)
g28358(1) = OR(g27149, g15837)
g33873(1) = AND(g33291, g20549)
g30033(1) = AND(g29189, g12937)
g28721(1) = OR(g27488, g16705)
g29523(1) = AND(g28930, g22417)
g29176(1) = OR(g27661, g17177)
g31292(1) = AND(g29735, g23338)
g29351(1) = AND(g4771, g28406)
g29516(1) = AND(g28895, g22369)
g32208(1) = OR(g31120, g29584)
g29208(1) = AND(g24138, I27538, I27539)
g31492(1) = AND(g29790, g23431)
g30029(1) = AND(g29164, g12936)
g29614(1) = AND(g28860, g22369)
g30028(1) = AND(g29069, g9311)
g31750(1) = AND(g30103, g23925)
g29607(1) = AND(g28509, g14208)
g29068(1) = OR(g27628, g17119)
g29593(1) = AND(g28470, g7985)
g29346(1) = AND(g4894, g28381)
g29565(1) = AND(g1932, g28590)
g29641(1) = AND(g28520, g14237)
g28347(1) = OR(g27138, g15822)
g29635(1) = AND(g28910, g22432)
g28420(1) = OR(g27222, g13290)
g29575(1) = AND(g2066, g28604)
g29327(1) = AND(g29070, g22156)
g28647(1) = OR(g27389, g16596)
g29537(1) = AND(g28976, g22472)
g29606(1) = AND(g28480, g8011)
g28296(1) = OR(g27095, g15784)
g28735(1) = OR(g27510, g16737)
g30045(1) = AND(g29200, g12419)
g31508(1) = AND(g29813, g23459)
g28345(1) = OR(g27137, g15821)
g28745(1) = OR(g27519, g16760)
g28814(1) = OR(g27545, g16841)
g30032(1) = AND(g29072, g9326)
g28600(1) = OR(g27339, g16427)
g29522(1) = AND(g28923, g22369)
g31756(1) = AND(g30114, g23942)
g29105(1) = OR(g27645, g17134)
g31780(1) = AND(g30163, g23999)
g29536(1) = AND(g28969, g22432)
g28305(1) = OR(g27103, g15793)
g32235(1) = OR(g31151, g29662)
g28699(1) = OR(g27452, g16667)
g28734(1) = OR(g27508, g16736)
g30071(1) = AND(g29184, g12975)
g34071(1) = AND(g8854, g33799)
g28556(1) = AND(g27431, g20374)
g32316(1) = AND(g31307, g23522)
g28401(1) = OR(g27212, g15871)
g29205(1) = AND(g24117, I27523, I27524)
g32247(1) = OR(g31168, g29686)
g28708(1) = OR(g27462, g16674)
g31769(1) = AND(g30141, g23986)
g29592(1) = AND(g28469, g11832)
g30059(1) = AND(g28106, g12467)
g30025(1) = AND(g28492, g23502)
g30058(1) = AND(g29180, g12950)
g29350(1) = AND(g4939, g28395)
g28668(1) = OR(g27411, g16617)
g30044(1) = AND(g29174, g12944)
g28850(1) = OR(g27557, g16869)
g33788(1) = OR(g33122, g32041)
g33710(1) = AND(g14037, g33246)
g31786(1) = AND(g30189, g24010)
g28293(1) = AND(g7424, g2495, g27474)
g32245(1) = OR(g31167, g29684)
g28334(1) = OR(g27131, g15817)
g28707(1) = OR(g27461, g16673)
g28206(1) = NAND(g12546, g26105, g27985)
g29640(1) = AND(g28498, g8125)
g28319(1) = OR(g27115, g15807)
g32216(1) = OR(g31128, g29615)
g29803(1) = AND(g28414, g26836)
g33717(1) = AND(g14092, g33306)
g28636(1) = OR(g27376, g16538)
g28419(1) = OR(g27221, g15884)
g29552(1) = AND(g2223, g28579)
g29204(1) = AND(g24110, I27518, I27519)
g28646(1) = OR(g27388, g16595)
g32227(1) = OR(g31146, g29648)
g28685(1) = OR(g27433, g16637)
g29647(1) = AND(g28934, g22457)
g28497(1) = OR(g27267, g16199)
g32277(1) = OR(g31211, g29733)
g32275(1) = OR(g31210, g29732)
g28744(1) = OR(g27518, g16759)
g29143(1) = OR(g27650, g17146)
g32308(1) = AND(g31293, g23503)
g30060(1) = AND(g29146, g10581)
g28661(1) = OR(g27406, g16611)
g28264(1) = AND(g7315, g1802, g27416)
g28667(1) = OR(g27410, g16616)
g28750(1) = OR(g27525, g16765)
g31765(1) = AND(g30128, g23968)
g29369(1) = AND(g28209, g22341)
g30070(1) = AND(g29167, g9529)
g33733(1) = OR(g33105, g32012)
g28542(1) = AND(g27405, g20275)
g31504(1) = AND(g29370, g10553)
g28453(1) = AND(g27582, g10233)
g29850(1) = AND(g28340, g24893)
g28530(1) = AND(g27383, g20240)
g28659(1) = OR(g27404, g16610)
g29627(1) = AND(g28493, g11884)
g29959(1) = AND(g28953, g12823)
g28288(1) = NAND(g10533, g26105, g27004)
g28490(1) = OR(g27262, g16185)
g32160(1) = AND(g31001, g22995)
g28749(1) = OR(g27523, g16764)
g28386(1) = OR(g27202, g13277)
g34157(1) = AND(g33794, g20159)
g31499(1) = AND(g29801, g23446)
g29548(1) = AND(g1798, g28575)
g28718(1) = OR(g27483, g16702)
g28283(1) = AND(g7380, g2361, g27445)
g28303(1) = AND(g7462, g2629, g27494)
g29626(1) = AND(g28584, g11415)
g32226(1) = OR(g31145, g29645)
g29533(1) = AND(g28958, g22417)
g32211(1) = OR(g31124, g29603)
g30596(1) = AND(g30279, g18947)
g28731(1) = OR(g27504, g16733)
g31132(1) = AND(g29504, g22987)
g28385(1) = OR(g27201, g15857)
g28778(1) = OR(g27540, g16808)
g28777(1) = OR(g27539, g16807)
g28635(1) = OR(g27375, g16537)
g31471(1) = AND(g29754, g23399)
g28252(1) = AND(g27159, g19682)
g29989(1) = AND(g29006, g10489)
g29611(1) = AND(g28540, g14209)
g29988(1) = AND(g29187, g12235)
g28684(1) = OR(g27432, g16636)
g28818(1) = OR(g27549, g13998)
g31792(1) = AND(g30214, g24017)
g32166(1) = AND(g31007, g23029)
g29650(1) = AND(g28949, g22472)
g28522(1) = NAND(g10857, g26131, g27142)
g28417(1) = OR(g27219, g15881)
g28373(1) = OR(g27180, g15849)
g28643(1) = OR(g27386, g16592)
g28623(1) = OR(g27361, g16520)
g31125(1) = AND(g29502, g22973)
g30015(1) = AND(g29040, g10519)
g28846(3) = AND(g21434, g26424, g25399, g27474)
g28259(1) = NAND(g10504, g26987, g26973)
g28287(1) = NAND(g10504, g26131, g26973)
g28702(1) = OR(g27457, g16670)
g29166(1) = OR(g27653, g17153)
g34084(1) = AND(g9214, g33851)
g31017(1) = AND(g29479, g22841)
g33732(1) = OR(g33104, g32011)
g32264(1) = OR(g31187, g29711)
g28634(1) = OR(g27374, g16536)
g28632(1) = OR(g27373, g16535)
g28641(1) = OR(g27385, g16591)
g29598(1) = AND(g28823, g22342)
g28691(1) = OR(g27437, g16642)
g28768(3) = AND(g21434, g26424, g25308, g27421)
g31752(1) = AND(g30104, g23928)
g31374(1) = AND(g29748, g23390)
g28429(1) = OR(g27228, g15913)
g28329(1) = OR(g27128, g15813)
g29656(1) = AND(g28515, g11666)
g29336(1) = AND(g4704, g28363)
g28730(1) = OR(g27503, g13912)
g31525(1) = AND(g29892, g23526)
g31016(1) = AND(g29478, g22840)
g28249(1) = AND(g27152, g19677)
g28717(1) = OR(g27482, g16701)
g29571(1) = AND(g28452, g11762)
g31270(1) = AND(g29692, g23282)
g30007(1) = AND(g29141, g12929)
g28516(1) = NAND(g10857, g26105, g27155)
g28511(1) = OR(g27272, g16208)
g28816(1) = OR(g27547, g16843)
g28372(1) = OR(g27178, g15848)
g31470(1) = AND(g29753, g23398)
g31494(1) = AND(g29792, g23435)
g28650(1) = OR(g27391, g16598)
g29610(1) = AND(g28483, g8026)
g28619(1) = OR(g27358, g16517)
g32237(1) = OR(g31153, g29667)
g30006(1) = AND(g29032, g9259)
g28701(1) = OR(g27455, g16669)
g28228(1) = AND(g27126, g19636)
g28746(1) = OR(g27520, g16762)
g28403(1) = OR(g27214, g13282)
g31477(1) = AND(g29763, g23409)
g28724(1) = OR(g27491, g16707)
g31118(1) = AND(g29490, g22906)
g28629(1) = OR(g27371, g16532)
g28774(1) = OR(g27536, g16804)
g31305(1) = AND(g29741, g23354)
g29201(1) = AND(g24081, I27503, I27504)
g28682(1) = OR(g27430, g16635)
g29595(1) = AND(g28475, g11833)
g28681(1) = OR(g27428, g16634)
g29623(1) = AND(g28496, g11563)
g28328(1) = OR(g27127, g15812)
g29352(1) = AND(g4950, g28410)
g28815(1) = OR(g27546, g16842)
g31485(1) = AND(g29776, g23421)
g30034(1) = AND(g29077, g10541)
g29836(1) = AND(g28425, g26841)
g28610(1) = OR(g27347, g16484)
g28295(1) = OR(g27094, g15783)
g28618(1) = OR(g27357, g16516)
g31519(1) = AND(g29864, g23490)
g28362(1) = OR(g27154, g15840)
g28880(3) = AND(g21434, g26424, g25438, g27494)
g28361(1) = OR(g27153, g15839)
g28851(1) = OR(g27558, g16870)
g28402(1) = OR(g27213, g15873)
g28207(1) = NAND(g12546, g26131, g27977)
g28628(1) = OR(g27370, g16531)
g32233(1) = OR(g31150, g29661)
g29555(1) = AND(g29004, g22498)
g28649(1) = OR(g27390, g16597)
g29567(1) = AND(g2357, g28593)
g29594(1) = AND(g28529, g14192)
g28172(1) = OR(g27469, g27440, g27416, g27395)
g32218(1) = OR(g31130, g29619)
g29518(1) = AND(g28906, g22384)
g31484(1) = AND(g29775, g23418)
g31115(1) = AND(g29487, g22882)
g29349(1) = AND(g4760, g28391)
g28688(1) = OR(g27435, g16639)
g33805(1) = AND(g33232, g20079)
g30047(1) = AND(g29109, g9407)
g28671(1) = OR(g27413, g16619)
g30592(1) = AND(g30270, g18929)
g32210(1) = OR(g31123, g29600)
g32209(1) = OR(g31122, g29599)
g28609(1) = OR(g27346, g16483)
g29554(1) = AND(g28997, g22472)
g29609(1) = AND(g28482, g11861)
g29608(1) = AND(g28568, g11385)
g28271(1) = NAND(g10533, g27004, g26990)
g29355(2) = NAND(g24383, g28109)
g28348(1) = OR(g27139, g15823)
g30046(1) = AND(g29108, g10564)
g29973(1) = AND(g28981, g9206)
g28357(1) = OR(g27148, g15836)
g32162(1) = AND(g31002, g23014)
g28571(1) = AND(g27458, g20435)
g28310(1) = OR(g27107, g15797)
g33759(1) = AND(g33123, g22847)
g29207(1) = AND(g24131, I27533, I27534)
g31758(1) = AND(g30115, g23945)
g31744(1) = AND(g30092, g23902)
g32229(1) = OR(g31148, g29652)
g30027(1) = AND(g29104, g12550)
I26741(1) = OR(g22881, g22905, g22928, g27402)
I29297(1) = NAND(g12117, I29295)
I26460(1) = NAND(g26576, I26459)
I29296(1) = NAND(g29495, I29295)
I26419(1) = NAND(g14247, I26417)
I26418(1) = NAND(g26519, I26417)
I29315(1) = NAND(g12154, I29313)
I29262(1) = NAND(g29485, I29261)
I29263(1) = NAND(g12046, I29261)
I26439(1) = NAND(g26549, I26438)
I29314(1) = NAND(g29501, I29313)
I29279(1) = NAND(g12081, I29277)
I29278(1) = NAND(g29488, I29277)
I29286(1) = NAND(g12085, I29284)
I29270(1) = NAND(g29486, I29269)
I29271(1) = NAND(g12050, I29269)
I26071(1) = NAND(g26026, I26070)
I26072(1) = NAND(g13517, I26070)
I26440(1) = NAND(g14271, I26438)
g29335(1) = NAND(g25540, g28131)
I26395(1) = NAND(g14227, I26393)
I26050(1) = NAND(g25997, I26049)
I26051(1) = NAND(g13500, I26049)
I29303(1) = NAND(g29496, I29302)
I26461(1) = NAND(g14306, I26459)
I26367(1) = NAND(g26400, I26366)
I26394(1) = NAND(g26488, I26393)
I26095(1) = NAND(g13539, I26093)
I26094(1) = NAND(g26055, I26093)
g29497(1) = NOR(g22763, g28241)
I29255(1) = NAND(g12017, I29253)
I29285(1) = NAND(g29489, I29284)
I26368(1) = NAND(g14211, I26366)
I29254(1) = NAND(g29482, I29253)
I29304(1) = NAND(g12121, I29302)
g29503(1) = NOR(g22763, g28250)
g31521(1) = NOT(I29182)
g33046(1) = OR(g32308, g21912)
g31877(1) = OR(g31278, g21732)
g30393(1) = OR(g29986, g21748)
g31880(1) = OR(g31280, g21774)
g31920(1) = OR(g31493, g22045)
g31925(1) = OR(g31789, g22061)
g29263(1) = OR(g28239, g18617)
g31869(1) = OR(g30592, g18221)
g33965(1) = OR(g33805, g18179)
g31924(1) = OR(g31486, g22049)
g30457(1) = OR(g29369, g21885)
g30414(1) = OR(g30002, g21794)
g31923(1) = OR(g31763, g22048)
g31882(1) = OR(g31115, g21776)
g29298(1) = OR(g28571, g18793)
g31878(1) = OR(g31015, g21733)
g31905(1) = OR(g31746, g21952)
g31886(1) = OR(g31481, g21791)
g31926(1) = OR(g31765, g22090)
g30480(1) = OR(g29321, g21972)
g31915(1) = OR(g31520, g22001)
g31917(1) = OR(g31478, g22003)
g33960(1) = OR(g33759, g21701)
g31890(1) = OR(g31143, g21823)
g31892(1) = OR(g31019, g21825)
g31899(1) = OR(g31470, g21907)
g31916(1) = OR(g31756, g22002)
g30459(1) = OR(g29314, g21926)
g30543(1) = OR(g29338, g22110)
g31912(1) = OR(g31752, g21998)
g31902(1) = OR(g31744, g21910)
g34022(1) = OR(g33873, g18538)
g29292(1) = OR(g28556, g18776)
g31891(1) = OR(g31305, g21824)
g31903(1) = OR(g31374, g21911)
g31887(1) = OR(g31292, g21820)
g31907(1) = OR(g31492, g21954)
g31875(1) = OR(g31066, g21730)
g29269(1) = OR(g28249, g18634)
g31909(1) = OR(g31750, g21956)
g31883(1) = OR(g31132, g21777)
g31874(1) = OR(g31016, g21729)
g33020(1) = OR(g32160, g21734)
g31910(1) = OR(g31471, g21957)
g31906(1) = OR(g31477, g21953)
g31918(1) = OR(g31786, g22015)
g31900(1) = OR(g31484, g21908)
g29304(1) = OR(g28588, g18810)
g33961(1) = OR(g33789, g21712)
g33025(1) = OR(g32162, g21780)
g31921(1) = OR(g31508, g22046)
g31879(1) = OR(g31475, g21745)
g30501(1) = OR(g29327, g22018)
g31893(1) = OR(g31490, g21837)
g31884(1) = OR(g31290, g21778)
g30435(1) = OR(g30025, g21840)
g31908(1) = OR(g31519, g21955)
g31876(1) = OR(g31125, g21731)
g31927(1) = OR(g31500, g22091)
g31919(1) = OR(g31758, g22044)
g31932(1) = OR(g31792, g22107)
g30522(1) = OR(g29332, g22064)
g31929(1) = OR(g31540, g22093)
g34251(1) = OR(g34157, g18147)
g31873(1) = OR(g31270, g21728)
g33061(1) = OR(g32334, g22050)
g31914(1) = OR(g31499, g22000)
g31930(1) = OR(g31769, g22094)
g29286(1) = OR(g28542, g18759)
g31889(1) = OR(g31118, g21822)
g31928(1) = OR(g31517, g22092)
g31911(1) = OR(g31784, g21969)
g31931(1) = OR(g31494, g22095)
g31881(1) = OR(g31018, g21775)
g31904(1) = OR(g31780, g21923)
g31871(1) = OR(g30596, g18279)
g33051(1) = OR(g32316, g21958)
g31913(1) = OR(g31485, g21999)
g33066(1) = OR(g32341, g22096)
g33056(1) = OR(g32327, g22004)
g31888(1) = OR(g31067, g21821)
g29222(1) = OR(g28252, g18105)
g31922(1) = OR(g31525, g22047)
g31901(1) = OR(g31516, g21909)
g33030(1) = OR(g32166, g21826)
g31898(1) = OR(g31707, g21906)
g29280(1) = OR(g28530, g18742)
g29257(1) = OR(g28228, g18600)
g31885(1) = OR(g31017, g21779)
g30326(1) = NOT(I28579)
g28367(1) = NOT(I26880)
g33250(1) = NOT(g32186)
g30614(55) = AND(g20154, g29814)
g30999(1) = NOT(g29722)
g30998(1) = NOT(g29719)
I28419(1) = NOT(g29195)
g30673(55) = AND(g20175, g29814)
g31672(33) = AND(g29814, g19050)
g30735(88) = AND(g29814, g22319)
g31376(88) = AND(g24952, g29814)
g30825(88) = AND(g29814, g22332)
g31528(11) = AND(g19050, g29814)
I28585(1) = NOT(g30217)
g28349(2) = NAND(g27074, g24770, g27187, g19644)
g31070(44) = AND(g29814, g25985)
g31194(11) = AND(g19128, g29814)
I26664(1) = NOT(g27708)
g30937(44) = AND(g22626, g29814)
g31170(11) = AND(g19128, g29814)
g31579(11) = AND(g19128, g29814)
I26687(1) = NOT(g27880)
g31710(33) = AND(g29814, g19128)
g31021(44) = AND(g26025, g29814)
I26705(1) = NOT(g27967)
I26679(1) = NOT(g27773)
g31154(11) = AND(g19128, g29814)
g29755(1) = NOT(I28002)
g30989(1) = NOT(g29672)
g28463(2) = NOT(I26952)
I26693(1) = NOT(g27930)
g30934(1) = NOR(g29836, g29850)
g29318(1) = NOT(g29029)
g30309(1) = NOT(g28959)
g32017(1) = NOR(g31504, g23475)
g31554(11) = AND(g19050, g29814)
g28752(1) = NOT(I27232)
g30195(1) = NOT(I28434)
g31327(44) = AND(g19200, g29814)
g28954(1) = NOT(g27830)
I29363(1) = NOT(g30218)
g29042(1) = NOT(I27388)
I27271(1) = NOT(g27998)
I26682(1) = NOT(g27774)
g30305(1) = NOT(g28939)
g31542(11) = AND(g19050, g29814)
I29204(1) = NOT(g29505)
g30565(1) = NOT(I28832)
I26785(1) = NOT(g27013)
g31667(1) = NOT(g30142)
g30567(1) = NOT(g29930)
g28224(1) = AND(g27163, g22763, g27064)
g30312(1) = NOT(g28970)
I26649(1) = NOT(g27675)
g31000(1) = NOT(g29737)
I28480(1) = NOT(g28652)
g31638(1) = NOT(g29689)
I26700(1) = NOT(g27956)
g28917(1) = NOT(I27314)
g28436(2) = NOT(I26929)
I27385(1) = NOT(g27438)
g31003(3) = NAND(g27163, g29497, g19644)
I27738(1) = NOT(g28140)
g31566(11) = AND(g19050, g29814)
I26670(1) = NOT(g27709)
g31522(1) = NOT(I29185)
g30990(1) = NOT(g29676)
g29384(1) = AND(g26424, g22763, g28179)
I29013(1) = NOT(g29705)
g30997(1) = NOT(g29702)
g30321(1) = NOT(I28572)
g30591(1) = NOT(I28851)
g34147(1) = NOT(g33823)
g30996(1) = NOT(g29694)
g29311(1) = NOT(g28998)
I29002(1) = NOT(g29675)
g30572(1) = NOT(g29945)
g30296(1) = NOT(g28889)
I26676(1) = NOT(g27736)
g28231(1) = AND(g27187, g22763, g27074)
I29337(1) = NOT(g30286)
g29043(1) = NOT(I27391)
g29310(1) = NOT(g28991)
g29765(1) = NOT(I28014)
g28336(2) = NAND(g27064, g24756, g27163, g19644)
g31008(1) = NOR(g30004, g30026)
I27481(1) = NOT(g27928)
g29013(1) = NOT(I27368)
g29365(1) = NOT(g29067)
g34359(3) = NOR(g9162, g34174, g12259)
g30568(1) = NOT(g29339)
g28779(1) = NOT(I27253)
g30578(1) = NOT(g29956)
g30983(1) = NOT(g29657)
g29382(1) = AND(g26424, g22763, g28172)
g31623(1) = NOT(g29669)
I28336(1) = NOT(g29147)
g34351(1) = NOT(g34174)
g30593(1) = NOT(g29970)
g34162(3) = NAND(g785, g33823, g11679)
g30929(1) = NOR(g29803, g29835)
g31653(1) = NOT(g29713)
g31608(1) = NOT(g29653)
g31009(3) = NAND(g27187, g29503, g19644)
g30302(1) = NOT(g28924)
g30248(1) = AND(g28743, g23938)
g29771(1) = AND(g28322, g23242)
g30204(1) = AND(g28670, g23868)
g33332(1) = AND(g32217, g20608)
g33361(1) = AND(g32257, g20911)
g30233(1) = AND(g28720, g23913)
g31257(1) = OR(g29531, g28253)
g31276(1) = OR(g29567, g28282)
g32120(1) = AND(g31639, g29941)
g32146(1) = AND(g31624, g29978)
g30143(1) = NOR(g28761, g14566)
g32408(1) = OR(g31541, g30073)
g29759(1) = AND(g28308, g23226)
g31267(1) = OR(g29548, g28263)
g29758(1) = AND(g28306, g23222)
g30212(1) = AND(g28687, g23879)
g31514(1) = AND(g20041, g29956)
g29962(1) = AND(g23616, g28959)
g32127(1) = AND(g31624, g29950)
g32103(1) = AND(g31609, g29905)
g33358(1) = AND(g32249, g20778)
g30229(1) = AND(g28716, g23904)
g33344(1) = AND(g32228, g20670)
g30228(1) = AND(g28715, g23903)
g29795(1) = AND(g28344, g23257)
g32126(1) = AND(g31601, g29948)
g29789(1) = AND(g28270, g10233)
g31466(1) = OR(g26160, g29650)
g29788(1) = AND(g28335, g23250)
g31990(1) = AND(g31772, g18945)
g30245(1) = AND(g28733, g23935)
g31306(1) = OR(g29595, g29610)
g29760(1) = AND(g28309, g23227)
g30232(1) = AND(g28719, g23912)
g32111(1) = AND(g31616, g29922)
g30261(1) = AND(g28772, g23961)
g30171(1) = NOR(g28880, g7431)
g30117(1) = NOR(g28739, g7252)
g32150(1) = AND(g31624, g29995)
g29199(1) = AND(g27187, g12687)
g29770(1) = AND(g28320, g23238)
g29767(1) = AND(g28317, g23236)
g29794(1) = AND(g28342, g23256)
g29845(1) = AND(g28375, g23291)
g29899(1) = AND(g28428, g23375)
g31249(1) = OR(g25971, g29523)
g30199(1) = AND(g28664, g23861)
g29718(1) = AND(g28512, g11136)
g30198(1) = AND(g28662, g23860)
g31274(1) = OR(g29565, g28280)
g32157(1) = AND(g31646, g30021)
g29861(1) = AND(g28390, g23313)
g33355(1) = AND(g32243, g20769)
g30225(1) = AND(g28705, g23897)
g31996(1) = AND(g31779, g18979)
g30258(1) = AND(g28751, g23953)
g33367(1) = AND(g32271, g21053)
g30244(1) = AND(g28732, g23930)
g28484(3) = AND(g27187, g10290, g21163, I26972)
g29766(1) = AND(g28316, g23235)
g34069(1) = AND(g8774, g33797)
g31304(1) = OR(g29594, g29608)
g29871(1) = AND(g28400, g23332)
g31291(1) = OR(g29581, g29593)
g31253(1) = OR(g25980, g29533)
g30106(1) = NOR(g28739, g7268)
g32156(1) = AND(g31639, g30018)
g30170(1) = NOR(g28846, g14615)
g29785(1) = AND(g28332, g23248)
g30599(1) = AND(g18911, g29863)
g30598(1) = AND(g18898, g29862)
g29859(1) = AND(g28388, g23307)
g29858(1) = AND(g28387, g23306)
g34322(1) = AND(g14188, g34174)
g29844(1) = AND(g28374, g23290)
g28539(1) = AND(g27187, g12762)
g32286(1) = AND(g31658, g29312)
g31289(1) = OR(g29580, g29591)
g27876(1) = NAND(I26418, I26419)
g32143(1) = AND(g31646, g29967)
g30144(1) = NOR(g28789, g7322)
g29902(1) = AND(g28430, g23377)
g30289(1) = AND(g28884, g24000)
g30224(1) = AND(g28704, g23896)
g29178(1) = AND(g27163, g12687)
g32110(1) = AND(g31639, g29921)
g31748(1) = NAND(I29303, I29304)
g31497(1) = AND(g20041, g29930)
g31747(1) = NAND(I29296, I29297)
g31767(1) = OR(g30031, g30043)
g28141(1) = AND(g10831, g11797, g11261, g27163)
g33339(1) = AND(g32221, g20634)
g30119(1) = NOR(g28761, g7315)
g33338(1) = AND(g32220, g20633)
g29784(1) = AND(g28331, g23247)
g31757(1) = OR(g29992, g30010)
g29888(1) = AND(g28418, g23352)
g30255(1) = AND(g28748, g23946)
g30188(1) = AND(g28644, g23841)
g31503(1) = AND(g20041, g29945)
g30267(1) = AND(g28776, g23967)
g31245(1) = OR(g25964, g29516)
g30219(1) = AND(g28698, g23887)
g29860(1) = AND(g28389, g23312)
g31766(1) = OR(g30029, g30042)
g29197(1) = OR(g27187, g27163)
g30277(1) = AND(g28817, g23987)
g30595(1) = AND(g18911, g29847)
g32116(1) = AND(g31658, g29929)
g30266(1) = AND(g28775, g23966)
g31468(1) = OR(g29641, g29656)
g29188(1) = AND(g27163, g12762)
g30148(1) = NOR(g28799, g7335)
g30167(1) = AND(g28622, g23793)
g30194(1) = AND(g28651, g23849)
g30589(1) = AND(g18898, g29811)
g32142(1) = AND(g31616, g29965)
g29979(1) = AND(g23655, g28991)
g31669(1) = NAND(I29254, I29255)
g29877(1) = AND(g28405, g23340)
g30254(1) = AND(g28747, g23944)
g30177(1) = AND(g28631, g23814)
g30183(1) = NOR(g28880, g14644)
g31709(1) = NAND(I29285, I29286)
g30166(1) = AND(g28621, g23792)
g33341(1) = AND(g32223, g20640)
g31774(1) = OR(g30046, g30057)
g30239(1) = AND(g28728, g23923)
g30594(1) = AND(g18898, g29846)
g29876(1) = AND(g28404, g23339)
g29885(1) = AND(g28416, g23350)
g30238(1) = AND(g28727, g23922)
g30185(1) = AND(g28640, g23838)
g30154(1) = AND(g28611, g23769)
g31256(1) = OR(g25983, g29537)
g30159(1) = NOR(g28799, g14589)
g32122(1) = AND(g31646, g29944)
g31269(1) = OR(g26024, g29569)
g32153(1) = AND(g31646, g29999)
g31761(1) = OR(g30009, g30028)
g30215(1) = AND(g28690, g23881)
g29773(1) = AND(g28203, g10233)
g27401(1) = NAND(I26094, I26095)
g30284(1) = AND(g28852, g23994)
g34348(1) = AND(g34125, g20128)
g33363(1) = AND(g32262, g20918)
g32109(1) = AND(g31609, g29920)
g32108(1) = AND(g31631, g29913)
g31223(1) = AND(g20028, g29689)
g31259(1) = OR(g25992, g29554)
g30146(1) = NOR(g28833, g7411)
g31708(1) = NAND(I29278, I29279)
g30576(1) = AND(g18898, g29800)
g30200(1) = AND(g28665, g23862)
g33334(1) = AND(g32219, g20613)
g31317(1) = OR(g29611, g29626)
g29373(1) = OR(g13832, g28453)
g29110(3) = AND(g27187, g12687, g20751, I27429)
g31760(1) = OR(g30007, g30027)
g30207(1) = AND(g28680, g23874)
g30005(1) = AND(g28230, g24394)
g31773(1) = OR(g30044, g30056)
g30241(1) = AND(g28729, g23926)
g31295(1) = OR(g26090, g29598)
g29762(1) = AND(g28298, g10233)
g30235(1) = AND(g28723, g23915)
g29909(1) = AND(g28435, g23388)
g30147(1) = NOR(g28768, g14567)
g29366(1) = OR(g13738, g28439)
g32152(1) = AND(g31631, g29998)
g29747(1) = AND(g28286, g23196)
g33340(1) = AND(g32222, g20639)
g29751(1) = AND(g28297, g23216)
g29807(1) = AND(g28359, g23272)
g29772(1) = AND(g28323, g23243)
g33362(1) = AND(g32259, g20914)
g29841(1) = AND(g28371, g23283)
g32113(1) = AND(g31601, g29925)
g31258(1) = OR(g25991, g29550)
g31279(1) = OR(g29571, g29579)
g30263(1) = AND(g28773, g23962)
g33351(1) = AND(g32236, g20707)
g33372(1) = AND(g32285, g21183)
g30221(1) = AND(g28700, g23893)
g29806(1) = AND(g28358, g23271)
g32248(1) = AND(g31616, g30299)
g30234(1) = AND(g28721, g23914)
g31753(1) = NAND(I29314, I29315)
g28150(1) = AND(g10862, g11834, g11283, g27187)
g29347(1) = AND(g29176, g22201)
g31322(1) = OR(g26128, g29635)
g29952(1) = AND(g23576, g28939)
g34107(1) = OR(g33710, g33121)
g32149(1) = AND(g31658, g29983)
g33327(1) = AND(g32208, g20561)
g32148(1) = AND(g31631, g29981)
g32104(1) = AND(g31616, g29906)
g31473(1) = OR(g26180, g29666)
g30156(1) = NOR(g28789, g14587)
g29320(1) = AND(g29068, g22147)
g29073(3) = AND(g27163, g10290, g21012, I27409)
g29797(1) = AND(g28347, g23259)
g27824(1) = NAND(I26394, I26395)
g30604(1) = AND(g18911, g29878)
g32112(1) = AND(g31646, g29923)
g29891(1) = AND(g28420, g23356)
g32096(1) = AND(g31601, g29893)
g30191(1) = AND(g28647, g23843)
g29750(1) = AND(g28296, g23215)
g29982(1) = AND(g23656, g28998)
g30247(1) = AND(g28735, g23937)
g29796(1) = AND(g28345, g23258)
g34324(1) = AND(g14064, g34161)
g30251(1) = AND(g28745, g23940)
g30272(1) = AND(g28814, g23982)
g32129(1) = AND(g31658, g29955)
g32128(1) = AND(g31631, g29953)
g29192(1) = AND(g27163, g10290)
g30140(1) = AND(g28600, g23749)
g31311(1) = OR(g26103, g29618)
g29949(1) = AND(g23575, g28924)
g31241(1) = OR(g25959, g29510)
g29326(1) = AND(g29105, g22155)
g29757(1) = AND(g28305, g23221)
g33350(1) = AND(g32235, g20702)
g31251(1) = OR(g25973, g29527)
g30220(1) = AND(g28699, g23888)
g30246(1) = AND(g28734, g23936)
g29872(1) = AND(g28401, g23333)
g30130(1) = NOR(g28761, g7275)
g32145(1) = AND(g31609, g29977)
g33357(1) = AND(g32247, g20775)
g30227(1) = AND(g28708, g23899)
g31320(1) = OR(g26125, g29632)
g30203(1) = AND(g28668, g23864)
g30281(1) = AND(g28850, g23992)
g32258(1) = AND(g31624, g30303)
g34146(1) = AND(g33788, g20091)
g32244(1) = AND(g31609, g30297)
g27767(1) = NAND(I26367, I26368)
g31465(1) = OR(g26156, g29647)
g33356(1) = AND(g32245, g20772)
g31706(1) = NAND(I29270, I29271)
g29787(1) = AND(g28334, g23249)
g30226(1) = AND(g28707, g23898)
g29743(1) = AND(g28206, g10233)
g29769(1) = AND(g28319, g23237)
g33331(1) = AND(g32216, g20607)
g31785(1) = OR(g30071, g30082)
g31751(1) = OR(g29975, g29990)
g31212(1) = AND(g20028, g29669)
g30181(1) = AND(g28636, g23821)
g31308(1) = OR(g26101, g29614)
g32159(1) = AND(g31658, g30040)
g29890(1) = AND(g28419, g23355)
g32158(1) = AND(g31658, g30022)
g30190(1) = AND(g28646, g23842)
g33343(1) = AND(g32227, g20665)
g30211(1) = AND(g28685, g23878)
g30024(1) = AND(g28497, g23501)
g33369(1) = AND(g32277, g21060)
g33368(1) = AND(g32275, g21057)
g29182(1) = AND(g27163, g12730)
g30250(1) = AND(g28744, g23939)
g31228(1) = AND(g20028, g29713)
g29331(1) = AND(g29143, g22169)
g27925(1) = NAND(I26439, I26440)
g30157(1) = NOR(g28833, g7369)
g30197(1) = AND(g28661, g23859)
g31745(1) = OR(g29959, g29973)
g31250(1) = OR(g25972, g29526)
g30202(1) = AND(g28667, g23863)
g30257(1) = AND(g28750, g23952)
g34111(1) = AND(g33733, g22936)
g30590(1) = AND(g18911, g29812)
g31248(1) = OR(g25970, g29522)
g31254(1) = OR(g25981, g29534)
g30196(1) = AND(g28659, g23858)
g30150(1) = NOR(g28846, g7424)
g30123(1) = NOR(g28768, g7328)
g30169(1) = NOR(g28833, g14613)
g29742(1) = AND(g28288, g10233)
g30001(1) = AND(g28490, g23486)
g30256(1) = AND(g28749, g23947)
g29857(1) = AND(g28386, g23304)
g27365(1) = NAND(I26050, I26051)
g30231(1) = AND(g28718, g23907)
g31770(1) = OR(g30034, g30047)
g31768(1) = OR(g30033, g30045)
g28982(3) = AND(g27163, g12687, g20682, I27349)
g31671(1) = NAND(I29262, I29263)
g33342(1) = AND(g32226, g20660)
g33330(1) = AND(g32211, g20588)
g32119(1) = AND(g31609, g29939)
g30243(1) = AND(g28731, g23929)
g31749(1) = OR(g29974, g29988)
g29856(1) = AND(g28385, g23303)
g30269(1) = AND(g28778, g23970)
g28553(1) = AND(g27187, g10290)
g31303(1) = OR(g29592, g29606)
g30268(1) = AND(g28777, g23969)
g32276(1) = AND(g31646, g30313)
g30180(1) = AND(g28635, g23820)
g31287(1) = OR(g29578, g28292)
g28528(1) = AND(g27187, g12730)
g30210(1) = AND(g28684, g23877)
g30278(1) = AND(g28818, g23988)
g31782(1) = OR(g30060, g30070)
g31755(1) = OR(g29991, g30008)
g31775(1) = OR(g30048, g30059)
g31781(1) = OR(g30058, g30069)
g29736(1) = AND(g28522, g10233)
g29887(1) = AND(g28417, g23351)
g29843(1) = AND(g28373, g23289)
g30187(1) = AND(g28643, g23840)
g30168(1) = AND(g28623, g23794)
g31764(1) = OR(g30015, g30032)
g29810(1) = AND(g28259, g11317)
g29774(1) = AND(g28287, g10233)
g30223(1) = AND(g28702, g23895)
g31754(1) = OR(g29989, g30006)
g29337(1) = AND(g29166, g22180)
g34110(1) = AND(g33732, g22935)
g33364(1) = AND(g32264, g20921)
g30179(1) = AND(g28634, g23819)
g30178(1) = AND(g28632, g23815)
g30186(1) = AND(g28641, g23839)
g30132(1) = NOR(g28789, g7362)
g31260(1) = OR(g25993, g29555)
g31284(1) = OR(g29575, g28290)
g32139(1) = AND(g31601, g29960)
g31762(1) = OR(g30011, g30030)
g30216(1) = AND(g28691, g23882)
g29901(1) = AND(g28429, g23376)
g31326(1) = OR(g29627, g29640)
g29783(1) = AND(g28329, g23246)
g30000(1) = AND(g23685, g29029)
g30242(1) = AND(g28730, g23927)
g29966(1) = AND(g23617, g28970)
g31302(1) = OR(g29590, g28302)
g32115(1) = AND(g31631, g29928)
g30230(1) = AND(g28717, g23906)
g31188(1) = AND(g20028, g29653)
g29752(1) = AND(g28516, g10233)
g30041(1) = AND(g28511, g23518)
g30275(1) = AND(g28816, g23984)
g29842(1) = AND(g28372, g23284)
g31244(1) = OR(g25963, g29515)
g30162(1) = NOR(g28880, g7462)
g27380(1) = NAND(I26071, I26072)
g30193(1) = AND(g28650, g23848)
g30165(1) = AND(g28619, g23788)
g33352(1) = AND(g32237, g20712)
g30129(1) = NOR(g28739, g14537)
g30222(1) = AND(g28701, g23894)
g29938(1) = AND(g23552, g28889)
g30253(1) = AND(g28746, g23943)
g29875(1) = AND(g28403, g23337)
g30236(1) = AND(g28724, g23916)
g32114(1) = AND(g31624, g29927)
g30175(1) = AND(g28629, g23813)
g32107(1) = AND(g31624, g29912)
g30160(1) = NOR(g28846, g7387)
g30264(1) = AND(g28774, g23963)
g30134(1) = NOR(g28768, g7280)
g32141(1) = AND(g31639, g29963)
g30209(1) = AND(g28682, g23876)
g32398(1) = OR(g31526, g30061)
g30208(1) = AND(g28681, g23875)
g32263(1) = AND(g31631, g30306)
g31325(1) = OR(g29625, g29639)
g29782(1) = AND(g28328, g23245)
g34332(1) = OR(g34071, g33723)
g30274(1) = AND(g28815, g23983)
g34073(1) = AND(g8948, g33823)
g30153(1) = AND(g28610, g23768)
g31255(1) = OR(g25982, g29536)
g32106(1) = AND(g31601, g29911)
g29749(1) = AND(g28295, g23214)
g32234(1) = AND(g31601, g30292)
g30164(1) = AND(g28618, g23787)
g29809(1) = AND(g28362, g23274)
g31518(1) = AND(g20041, g29970)
g29808(1) = AND(g28361, g23273)
g29036(3) = AND(g27163, g12762, g20875, I27381)
g30283(1) = AND(g28851, g23993)
g29874(1) = AND(g28402, g23336)
g29693(1) = AND(g28207, g10233)
g31316(1) = OR(g29609, g29624)
g27955(1) = NAND(I26460, I26461)
g30174(1) = AND(g28628, g23812)
g29008(3) = AND(g27163, g12730, g20739, I27364)
g33349(1) = AND(g32233, g20699)
g32121(1) = AND(g31616, g29942)
g30192(1) = AND(g28649, g23847)
g31268(1) = OR(g29552, g28266)
g33333(1) = AND(g32218, g20612)
g28471(3) = AND(g27187, g12762, g21024, I26960)
g30136(1) = NOR(g28799, g7380)
g30213(1) = AND(g28688, g23880)
g30205(1) = AND(g28671, g23869)
g28458(3) = AND(g27187, g12730, g20887, I26948)
g33329(1) = AND(g32210, g20585)
g31315(1) = OR(g29607, g29623)
g33328(1) = AND(g32209, g20584)
g30152(1) = AND(g28609, g23767)
g32272(1) = AND(g31639, g30310)
g32140(1) = AND(g31609, g29961)
g29799(1) = AND(g28271, g10233)
g30583(5) = AND(g19666, g29355)
g29798(1) = AND(g28348, g23260)
g29805(1) = AND(g28357, g23270)
g29761(1) = AND(g28310, g23228)
g31246(1) = OR(g25965, g29518)
g32147(1) = AND(g31616, g29980)
g33345(1) = AND(g32229, g20671)
g32151(1) = AND(g31639, g29996)
I28566(1) = OR(g29201, g29202, g29203, g28035)
I28567(1) = OR(g29204, g29205, g29206, g29207)
g28220(2) = OR(g23495, I26741, I26742)
g29520(1) = OR(g28291, g28281, g28264, g28254)
g29529(1) = OR(g28303, g28293, g28283, g28267)
g30580(2) = NAND(g29335, g19666)
g30573(2) = NAND(g29355, g19666)
g33669(1) = NAND(g33378, g862)
g30405(1) = OR(g29767, g21764)
g30416(1) = OR(g29858, g21800)
g30466(1) = OR(g30174, g21937)
g30505(1) = OR(g30168, g22026)
g30432(1) = OR(g29888, g21816)
g33550(1) = OR(g33342, g18338)
g30494(1) = OR(g30209, g21990)
g34252(1) = OR(g34146, g18180)
g30489(1) = OR(g30250, g21985)
g30496(1) = OR(g30231, g21992)
g30533(1) = OR(g30203, g22079)
g30490(1) = OR(g30167, g21986)
g30427(1) = OR(g29796, g21811)
g33571(1) = OR(g33367, g18409)
g30534(1) = OR(g30213, g22080)
g30498(1) = OR(g30251, g21994)
g34438(1) = OR(g34348, g18150)
g30439(1) = OR(g29761, g21848)
g30541(1) = OR(g30281, g22087)
g30519(1) = OR(g30264, g22040)
g30476(1) = OR(g30229, g21947)
g30429(1) = OR(g29844, g21813)
g30424(1) = OR(g29760, g21808)
g30420(1) = OR(g29769, g21804)
g30404(1) = OR(g29758, g21763)
g30483(1) = OR(g30241, g21979)
g30453(1) = OR(g29902, g21862)
g30526(1) = OR(g30181, g22072)
g30499(1) = OR(g30261, g21995)
g30528(1) = OR(g30202, g22074)
g30521(1) = OR(g29331, g22042)
g30474(1) = OR(g30208, g21945)
g30510(1) = OR(g30263, g22031)
g33548(1) = OR(g33327, g18336)
g33588(1) = OR(g33334, g18468)
g30495(1) = OR(g30222, g21991)
g30403(1) = OR(g29750, g21762)
g30419(1) = OR(g29759, g21803)
g30504(1) = OR(g30253, g22025)
g30455(1) = OR(g30041, g21864)
g30444(1) = OR(g29901, g21853)
g30328(1) = NOT(I28585)
g30502(1) = OR(g30232, g22023)
g30555(1) = OR(g30227, g22126)
g30538(1) = OR(g30256, g22084)
g30497(1) = OR(g30242, g21993)
g30418(1) = OR(g29751, g21802)
g30438(1) = OR(g29890, g21847)
g30540(1) = OR(g30275, g22086)
g32986(1) = OR(g31996, g18280)
g30421(1) = OR(g29784, g21805)
g33573(1) = OR(g33343, g18415)
g30481(1) = OR(g30221, g21977)
g30517(1) = OR(g30244, g22038)
g30539(1) = OR(g30267, g22085)
g30436(1) = OR(g29860, g21845)
g30553(1) = OR(g30205, g22124)
g34250(1) = OR(g34111, g21713)
g32983(1) = OR(g31990, g18222)
g30402(1) = OR(g29871, g21761)
g30558(1) = OR(g30258, g22129)
g30462(1) = OR(g30228, g21933)
g30487(1) = OR(g30187, g21983)
g30531(1) = OR(g30274, g22077)
g30506(1) = OR(g30179, g22027)
g30451(1) = OR(g29877, g21860)
g30552(1) = OR(g30283, g22123)
g33595(1) = OR(g33368, g18489)
g33589(1) = OR(g33340, g18469)
g30557(1) = OR(g30247, g22128)
g30516(1) = OR(g30233, g22037)
g30486(1) = OR(g30177, g21982)
g30440(1) = OR(g29771, g21849)
g30530(1) = OR(g30224, g22076)
g30542(1) = OR(g29337, g22088)
g33597(1) = OR(g33344, g18495)
g30524(1) = OR(g30255, g22070)
g30475(1) = OR(g30220, g21946)
g30518(1) = OR(g30254, g22039)
g30450(1) = OR(g29861, g21859)
g34249(1) = OR(g34110, g21702)
g30523(1) = OR(g30245, g22069)
g30551(1) = OR(g30235, g22122)
g30452(1) = OR(g29891, g21861)
g30463(1) = OR(g30140, g21934)
g30546(1) = OR(g30277, g22117)
g30556(1) = OR(g30236, g22127)
g30428(1) = OR(g29807, g21812)
g30485(1) = OR(g30166, g21981)
g30422(1) = OR(g29795, g21806)
g30423(1) = OR(g29887, g21807)
g30529(1) = OR(g30212, g22075)
g33587(1) = OR(g33363, g18463)
g30460(1) = OR(g30207, g21931)
g30401(1) = OR(g29782, g21760)
g30411(1) = OR(g29872, g21770)
g33556(1) = OR(g33329, g18362)
g30472(1) = OR(g30186, g21943)
g30406(1) = OR(g29783, g21765)
g33603(1) = OR(g33372, g18515)
g33604(1) = OR(g33345, g18520)
g30415(1) = OR(g29843, g21799)
g30413(1) = OR(g30001, g21772)
g30549(1) = OR(g30215, g22120)
g30433(1) = OR(g29899, g21817)
g30478(1) = OR(g30248, g21949)
g33598(1) = OR(g33364, g18496)
g30468(1) = OR(g30238, g21939)
g30559(1) = OR(g30269, g22130)
g33557(1) = OR(g33331, g18363)
g30511(1) = OR(g30180, g22032)
g33563(1) = OR(g33361, g18383)
g33582(1) = OR(g33351, g18444)
g33581(1) = OR(g33333, g18443)
g30509(1) = OR(g30210, g22030)
g30445(1) = OR(g29772, g21854)
g30514(1) = OR(g30211, g22035)
g30493(1) = OR(g30198, g21989)
g30488(1) = OR(g30197, g21984)
g33580(1) = OR(g33330, g18442)
g30532(1) = OR(g30193, g22078)
g33564(1) = OR(g33332, g18388)
g30443(1) = OR(g29808, g21852)
g30508(1) = OR(g30199, g22029)
g30464(1) = OR(g30152, g21935)
g33606(1) = OR(g33369, g18522)
g30482(1) = OR(g30230, g21978)
g30525(1) = OR(g30266, g22071)
g30448(1) = OR(g29809, g21857)
g30513(1) = OR(g30200, g22034)
g30469(1) = OR(g30153, g21940)
g30548(1) = OR(g30204, g22119)
g30560(1) = OR(g30278, g22131)
g30431(1) = OR(g29875, g21815)
g30467(1) = OR(g30185, g21938)
g30442(1) = OR(g29797, g21851)
g30484(1) = OR(g30154, g21980)
g30527(1) = OR(g30192, g22073)
g30447(1) = OR(g29798, g21856)
g30562(1) = OR(g30289, g22133)
g30545(1) = OR(g30268, g22116)
g33590(1) = OR(g33358, g18470)
g30477(1) = OR(g30239, g21948)
g33579(1) = OR(g33357, g18437)
g30425(1) = OR(g29770, g21809)
g30507(1) = OR(g30190, g22028)
g33605(1) = OR(g33352, g18521)
g33558(1) = OR(g33350, g18364)
g30512(1) = OR(g30191, g22033)
g33572(1) = OR(g33339, g18414)
g30471(1) = OR(g30175, g21942)
g33555(1) = OR(g33355, g18357)
g30554(1) = OR(g30216, g22125)
g30537(1) = OR(g30246, g22083)
g30441(1) = OR(g29787, g21850)
g30446(1) = OR(g29788, g21855)
g30399(1) = OR(g29757, g21758)
g30547(1) = OR(g30194, g22118)
g30544(1) = OR(g30257, g22115)
g30561(1) = OR(g30284, g22132)
g30430(1) = OR(g29859, g21814)
g33565(1) = OR(g33338, g18389)
g33566(1) = OR(g33356, g18390)
g30465(1) = OR(g30164, g21936)
g30396(1) = OR(g29856, g21755)
g30520(1) = OR(g30272, g22041)
g30397(1) = OR(g29747, g21756)
g30409(1) = OR(g29842, g21768)
g30470(1) = OR(g30165, g21941)
g30398(1) = OR(g29749, g21757)
g30426(1) = OR(g29785, g21810)
g30515(1) = OR(g30223, g22036)
g30417(1) = OR(g29874, g21801)
g33574(1) = OR(g33362, g18416)
g30410(1) = OR(g29857, g21769)
g30454(1) = OR(g29909, g21863)
g33547(1) = OR(g33349, g18331)
g33596(1) = OR(g33341, g18494)
g33549(1) = OR(g33328, g18337)
g30408(1) = OR(g29806, g21767)
g30503(1) = OR(g30243, g22024)
g30550(1) = OR(g30226, g22121)
g30492(1) = OR(g30188, g21988)
g30536(1) = OR(g30234, g22082)
g30449(1) = OR(g29845, g21858)
g30461(1) = OR(g30219, g21932)
g30563(1) = OR(g29347, g22134)
g30437(1) = OR(g29876, g21846)
g30412(1) = OR(g29885, g21771)
g30491(1) = OR(g30178, g21987)
g30434(1) = OR(g30024, g21818)
g30479(1) = OR(g29320, g21950)
g30535(1) = OR(g30225, g22081)
g30394(1) = OR(g29805, g21753)
g30395(1) = OR(g29841, g21754)
g30458(1) = OR(g30005, g24330)
g30400(1) = OR(g29766, g21759)
g30473(1) = OR(g30196, g21944)
g30407(1) = OR(g29794, g21766)
g30500(1) = OR(g29326, g21996)
I28349(1) = NOT(g28367)
g30601(2) = NOR(g16279, g29718)
g33804(1) = NOT(g33250)
g31596(4) = NOT(I29204)
g32540(1) = NOT(g30614)
g30182(1) = NOT(I28419)
g32902(1) = NOT(g30673)
g32957(1) = NOT(g31672)
g30984(4) = OR(g29765, g29755)
g32739(1) = NOT(g30735)
g32738(1) = NOT(g31376)
g32562(1) = NOT(g30673)
g32645(1) = NOT(g30825)
g32699(1) = NOT(g31528)
g29725(4) = NOT(g28349)
g32698(1) = NOT(g30614)
g32632(1) = NOT(g31070)
g32661(1) = NOT(g31070)
g32547(1) = NOT(g30614)
g32895(1) = NOT(g30673)
g32481(1) = NOT(g31194)
g32551(1) = NOT(g30735)
g32572(1) = NOT(g30735)
g32490(1) = NOT(g30673)
g32784(1) = NOT(g31672)
g32956(1) = NOT(g30825)
g32889(1) = NOT(g31376)
g32888(1) = NOT(g30673)
g32824(1) = NOT(g31376)
g28155(1) = NOT(I26664)
g32671(1) = NOT(g31528)
g32931(1) = NOT(g30937)
I27735(1) = NOT(g28779)
g28166(1) = NOT(I26687)
g32546(1) = NOT(g31170)
I29582(1) = NOT(g30591)
g32860(1) = NOT(g30673)
g32497(1) = NOT(g30673)
g32700(1) = NOT(g31579)
g32659(1) = NOT(g30735)
g32625(1) = NOT(g31070)
g32658(1) = NOT(g31579)
g32943(1) = NOT(g31710)
g32644(1) = NOT(g30735)
g32969(1) = NOT(g30735)
g32968(1) = NOT(g31376)
I27718(1) = NOT(g28231)
g32855(1) = NOT(g30825)
g32870(1) = NOT(g31021)
g32527(1) = NOT(g30673)
I29368(1) = NOT(g30321)
g32503(1) = NOT(g31194)
g32867(1) = NOT(g30673)
g32894(1) = NOT(g30614)
g32581(1) = NOT(g31070)
g32714(1) = NOT(g31528)
g32707(1) = NOT(g31579)
g32819(1) = NOT(g30825)
g32818(1) = NOT(g30735)
g32496(1) = NOT(g30614)
g32590(1) = NOT(g31154)
g32741(1) = NOT(g31710)
g32801(1) = NOT(g30937)
g32735(1) = NOT(g31021)
g32877(1) = NOT(g30825)
I27777(1) = NOT(g29043)
g32695(1) = NOT(g30735)
g32526(1) = NOT(g30614)
g32457(1) = NOT(g30735)
g32866(1) = NOT(g30614)
g32917(1) = NOT(g30937)
g32706(1) = NOT(g30673)
g32597(1) = NOT(g31154)
g32689(1) = NOT(g30825)
g32923(1) = NOT(g31021)
g32688(1) = NOT(g30735)
g32624(1) = NOT(g30825)
g28162(1) = NOT(I26679)
g32876(1) = NOT(g30735)
g32885(1) = NOT(g31021)
g32854(1) = NOT(g30735)
g30259(1) = NOT(g28463)
g32511(1) = NOT(g30614)
g32763(1) = NOT(g31710)
g31771(1) = NOT(I29337)
g32660(1) = NOT(g30825)
g32456(1) = NOT(g31376)
g32480(1) = NOT(g31070)
g32916(1) = NOT(g31021)
g32550(1) = NOT(g31376)
g32721(1) = NOT(g31021)
g32596(1) = NOT(g31070)
g32773(1) = NOT(g31376)
g32942(1) = NOT(g30825)
g32655(1) = NOT(g30614)
g28184(1) = NOT(I26705)
g32670(1) = NOT(g30673)
g32734(1) = NOT(g31710)
g32839(1) = NOT(g30735)
g32930(1) = NOT(g31021)
g32667(1) = NOT(g30825)
g32694(1) = NOT(g31376)
g32838(1) = NOT(g31376)
g32965(1) = NOT(g31710)
g32487(1) = NOT(g30825)
g32619(1) = NOT(g30614)
g32502(1) = NOT(g31070)
g32557(1) = NOT(g31376)
g32618(1) = NOT(g31154)
g32469(1) = NOT(g30673)
I28540(1) = NOT(g28954)
g32468(1) = NOT(g30614)
g32038(1) = NOT(g30934)
g32815(1) = NOT(g30937)
g32601(1) = NOT(g31376)
g32677(1) = NOT(g30673)
g31950(8) = NAND(g7285, g30573)
g32937(1) = NOT(g31021)
g32329(1) = NOT(g31522)
g32791(1) = NOT(g31672)
g32884(1) = NOT(g30825)
g32479(1) = NOT(g30735)
g32666(1) = NOT(g31376)
g32478(1) = NOT(g31376)
g28819(1) = NOT(I27271)
g32486(1) = NOT(g30735)
g33426(1) = NOT(g32017)
g32556(1) = NOT(g31554)
g32580(1) = NOT(g30825)
I27730(1) = NOT(g28752)
g32922(1) = NOT(g31710)
g28161(1) = NOT(I26676)
g32531(1) = NOT(g31070)
g32740(1) = NOT(g31672)
g32676(1) = NOT(g30614)
g32685(1) = NOT(g31528)
g32953(1) = NOT(g31327)
g32654(1) = NOT(g31070)
g32800(1) = NOT(g31021)
g32936(1) = NOT(g31710)
g31189(4) = NOT(I29002)
g32762(1) = NOT(g31672)
g32964(1) = NOT(g31672)
g32587(1) = NOT(g30735)
g32909(1) = NOT(g30614)
g32543(1) = NOT(g31376)
g32908(1) = NOT(g31327)
g32569(1) = NOT(g30673)
g32568(1) = NOT(g31170)
g32747(1) = NOT(g30825)
g32814(1) = NOT(g31021)
g32751(1) = NOT(g31327)
g32807(1) = NOT(g31021)
g32772(1) = NOT(g31327)
g32974(1) = NOT(g30937)
g32639(1) = NOT(g31070)
g32638(1) = NOT(g30825)
g32841(1) = NOT(g31672)
g32510(1) = NOT(g31194)
g32579(1) = NOT(g30735)
I28301(1) = NOT(g29042)
g32578(1) = NOT(g31376)
g32835(1) = NOT(g31710)
g28163(1) = NOT(I26682)
g32586(1) = NOT(g31376)
g31213(4) = NOT(I29013)
g32615(1) = NOT(g31376)
g32720(1) = NOT(g31710)
g32746(1) = NOT(g30735)
g32493(1) = NOT(g30735)
g32465(1) = NOT(g30825)
g32806(1) = NOT(g31710)
g32684(1) = NOT(g30673)
g28173(1) = NOT(I26693)
g32517(1) = NOT(g31194)
g32523(1) = NOT(g30825)
g31791(1) = NOT(I29363)
g32475(1) = NOT(g30614)
g32727(1) = NOT(g31710)
g32863(1) = NOT(g31021)
g32703(1) = NOT(g30825)
g32600(1) = NOT(g31542)
g32781(1) = NOT(g31376)
g32952(1) = NOT(g30937)
g32821(1) = NOT(g31021)
g32790(1) = NOT(g30825)
g32516(1) = NOT(g31070)
I29579(1) = NOT(g30565)
g28262(1) = NOT(I26785)
g32873(1) = NOT(g30614)
g32834(1) = NOT(g31672)
g32542(1) = NOT(g31554)
I29149(1) = NOT(g29384)
g32726(1) = NOT(g31672)
g32913(1) = NOT(g30825)
g32614(1) = NOT(g31542)
g32607(1) = NOT(g31542)
g32905(1) = NOT(g30825)
g32530(1) = NOT(g30825)
g32593(1) = NOT(g31542)
g32565(1) = NOT(g30735)
g32464(1) = NOT(g30735)
g32641(1) = NOT(g30614)
g32797(1) = NOT(g30825)
g32635(1) = NOT(g31542)
g32891(1) = NOT(g30825)
I29139(1) = NOT(g29382)
g32575(1) = NOT(g31170)
g32474(1) = NOT(g31194)
g32711(1) = NOT(g31070)
g32537(1) = NOT(g30825)
g32606(1) = NOT(g30673)
g32492(1) = NOT(g31376)
g32750(1) = NOT(g30937)
g29730(1) = OR(g28150, g28141)
g32796(1) = NOT(g31376)
I27713(1) = NOT(g28224)
g32840(1) = NOT(g30825)
g32522(1) = NOT(g30735)
g32663(1) = NOT(g30673)
g30605(1) = OR(g29529, g29520)
g32483(1) = NOT(g30673)
g32553(1) = NOT(g31170)
g32862(1) = NOT(g30825)
g32949(1) = NOT(g30825)
g32536(1) = NOT(g31376)
g32948(1) = NOT(g30735)
g32702(1) = NOT(g30735)
g32757(1) = NOT(g30937)
g32904(1) = NOT(g30735)
g32621(1) = NOT(g31542)
g32564(1) = NOT(g31376)
g32673(1) = NOT(g31376)
g32847(1) = NOT(g30735)
g32509(1) = NOT(g31070)
g32933(1) = NOT(g31376)
g32508(1) = NOT(g30825)
g32634(1) = NOT(g30673)
g32851(1) = NOT(g31327)
g32872(1) = NOT(g31327)
g34354(3) = NOR(g9003, g34162, g11083)
g32574(1) = NOT(g31070)
g32912(1) = NOT(g30735)
g29372(1) = NOT(I27738)
g32592(1) = NOT(g30673)
g32756(1) = NOT(g31021)
g32820(1) = NOT(g31672)
g28181(1) = NOT(I26700)
g32846(1) = NOT(g31376)
I27749(1) = NOT(g28917)
g32731(1) = NOT(g31376)
g32072(9) = NAND(g31009, g13301)
g30206(1) = NOT(g28436)
g32691(1) = NOT(g30673)
g32929(1) = NOT(g31710)
g32583(1) = NOT(g30614)
g32928(1) = NOT(g31672)
g32787(1) = NOT(g30937)
g32743(1) = NOT(g30937)
g32827(1) = NOT(g31672)
g32640(1) = NOT(g31154)
g32769(1) = NOT(g31672)
g28142(1) = NOT(I26649)
g32768(1) = NOT(g30825)
g32803(1) = NOT(g31376)
g29041(1) = NOT(I27385)
g32881(1) = NOT(g30673)
g32662(1) = NOT(g30614)
g32890(1) = NOT(g30735)
g32482(1) = NOT(g30614)
g32710(1) = NOT(g30825)
g32552(1) = NOT(g30825)
g32779(1) = NOT(g30937)
g32778(1) = NOT(g31021)
g32786(1) = NOT(g31021)
g32647(1) = NOT(g31154)
g32945(1) = NOT(g30937)
g32826(1) = NOT(g30825)
g32090(3) = NOT(g31003)
g32651(1) = NOT(g31376)
g32672(1) = NOT(g31579)
g32932(1) = NOT(g31327)
g32513(1) = NOT(g31376)
g32897(1) = NOT(g30735)
g32961(1) = NOT(g31376)
g32505(1) = NOT(g31566)
g32057(9) = NAND(g31003, g13297)
g32717(1) = NOT(g30735)
g32723(1) = NOT(g31327)
g32620(1) = NOT(g30673)
g32811(1) = NOT(g30735)
g32646(1) = NOT(g31070)
g28157(1) = NOT(I26670)
g32971(1) = NOT(g31672)
g32850(1) = NOT(g30937)
g32896(1) = NOT(g31376)
g32716(1) = NOT(g31376)
g32582(1) = NOT(g31170)
g32627(1) = NOT(g30673)
g32959(1) = NOT(g30937)
g32925(1) = NOT(g31327)
g32958(1) = NOT(g31710)
g32603(1) = NOT(g31070)
g32742(1) = NOT(g31021)
g32944(1) = NOT(g31021)
g32681(1) = NOT(g30735)
g32802(1) = NOT(g31327)
g32857(1) = NOT(g30937)
g32730(1) = NOT(g31327)
g32793(1) = NOT(g31021)
g32765(1) = NOT(g31327)
g32690(1) = NOT(g31070)
g32549(1) = NOT(g31554)
g32548(1) = NOT(g30673)
g32504(1) = NOT(g30673)
g32626(1) = NOT(g30614)
g32533(1) = NOT(g30614)
g32775(1) = NOT(g30825)
g32737(1) = NOT(g31327)
g32697(1) = NOT(g31070)
g32856(1) = NOT(g31021)
g32880(1) = NOT(g30614)
g32512(1) = NOT(g31566)
g31971(2) = NAND(g30573, g10511)
g32831(1) = NOT(g31376)
g32499(1) = NOT(g31376)
g32498(1) = NOT(g31566)
g32611(1) = NOT(g31154)
g32722(1) = NOT(g30937)
g32924(1) = NOT(g30937)
g32753(1) = NOT(g30735)
g32461(1) = NOT(g30614)
g32736(1) = NOT(g30937)
g32887(1) = NOT(g30614)
g32529(1) = NOT(g30735)
g32528(1) = NOT(g31554)
g32696(1) = NOT(g30825)
g32843(1) = NOT(g31021)
g30922(2) = NOR(g16662, g29810)
g32764(1) = NOT(g30937)
g32869(1) = NOT(g30735)
g32960(1) = NOT(g31327)
g32868(1) = NOT(g31376)
g32709(1) = NOT(g30735)
g32708(1) = NOT(g31376)
g32471(1) = NOT(g31376)
g29185(1) = NOT(I27481)
g34550(2) = NAND(g626, g34359, g12323)
g32602(1) = NOT(g30825)
g32810(1) = NOT(g31376)
g32657(1) = NOT(g31528)
g32774(1) = NOT(g30735)
g32955(1) = NOT(g30735)
g32879(1) = NOT(g31327)
g32970(1) = NOT(g30825)
g32878(1) = NOT(g30937)
g32886(1) = NOT(g31327)
g32792(1) = NOT(g31710)
g32967(1) = NOT(g31327)
g32459(1) = NOT(g31070)
g32919(1) = NOT(g30735)
g32458(1) = NOT(g30825)
g32918(1) = NOT(g31327)
g32545(1) = NOT(g31070)
g32599(1) = NOT(g30673)
g32598(1) = NOT(g30614)
g32817(1) = NOT(g31376)
g32532(1) = NOT(g31170)
g32901(1) = NOT(g31327)
g32783(1) = NOT(g30825)
g30237(1) = NOT(I28480)
g32561(1) = NOT(g30614)
g32656(1) = NOT(g30673)
g32680(1) = NOT(g31376)
g32823(1) = NOT(g31327)
g32966(1) = NOT(g31021)
g32631(1) = NOT(g30825)
g32571(1) = NOT(g31376)
g32495(1) = NOT(g31070)
g32816(1) = NOT(g31327)
g32687(1) = NOT(g31376)
g32752(1) = NOT(g31376)
g32954(1) = NOT(g31376)
g32643(1) = NOT(g31376)
g32669(1) = NOT(g30614)
g32668(1) = NOT(g31070)
g32842(1) = NOT(g31710)
g32489(1) = NOT(g30614)
g32559(1) = NOT(g30825)
g32525(1) = NOT(g31170)
g32488(1) = NOT(g31194)
g32558(1) = NOT(g30735)
g32830(1) = NOT(g31327)
g32893(1) = NOT(g30937)
g32544(1) = NOT(g30735)
g32865(1) = NOT(g31327)
g32713(1) = NOT(g30673)
g32610(1) = NOT(g31070)
g32705(1) = NOT(g30614)
g32679(1) = NOT(g31579)
g32678(1) = NOT(g31528)
g32460(1) = NOT(g31194)
g32686(1) = NOT(g31579)
g32939(1) = NOT(g31327)
g32938(1) = NOT(g30937)
g32875(1) = NOT(g31376)
g32837(1) = NOT(g31327)
g32617(1) = NOT(g30825)
g32470(1) = NOT(g31566)
g32915(1) = NOT(g31710)
g32595(1) = NOT(g30825)
g32467(1) = NOT(g31194)
g32494(1) = NOT(g30825)
g32623(1) = NOT(g30735)
g32782(1) = NOT(g30735)
g32822(1) = NOT(g30937)
g32853(1) = NOT(g30673)
g32589(1) = NOT(g31070)
g32588(1) = NOT(g30825)
g32524(1) = NOT(g31070)
g32836(1) = NOT(g31021)
g32477(1) = NOT(g31566)
g29697(4) = NOT(g28336)
g32118(1) = NOT(g31008)
g32864(1) = NOT(g30937)
g32749(1) = NOT(g31021)
g32616(1) = NOT(g30735)
g32748(1) = NOT(g31710)
g32704(1) = NOT(g31070)
I29939(1) = NOT(g31667)
g32809(1) = NOT(g31327)
g32900(1) = NOT(g30937)
g32466(1) = NOT(g31070)
g32808(1) = NOT(g30937)
g32560(1) = NOT(g31070)
I27784(1) = NOT(g29013)
g32642(1) = NOT(g31542)
g32733(1) = NOT(g31672)
g32874(1) = NOT(g30673)
g29987(1) = AND(g29197, g26424, g22763)
g32630(1) = NOT(g30735)
g32693(1) = NOT(g31579)
g32665(1) = NOT(g31579)
g32892(1) = NOT(g31021)
g32476(1) = NOT(g30673)
g32485(1) = NOT(g31376)
g32555(1) = NOT(g30673)
g32570(1) = NOT(g31554)
g32712(1) = NOT(g30614)
g32914(1) = NOT(g31672)
g32907(1) = NOT(g30937)
g32567(1) = NOT(g31070)
g32594(1) = NOT(g30735)
g32941(1) = NOT(g30735)
g32519(1) = NOT(g30673)
g32675(1) = NOT(g31070)
g32518(1) = NOT(g30614)
g32637(1) = NOT(g30735)
g32935(1) = NOT(g31672)
g32883(1) = NOT(g30735)
g32501(1) = NOT(g30825)
g32729(1) = NOT(g30937)
g32577(1) = NOT(g31554)
g32728(1) = NOT(g31021)
g32906(1) = NOT(g31021)
g32622(1) = NOT(g31376)
g32566(1) = NOT(g30825)
g32653(1) = NOT(g30825)
g32636(1) = NOT(g31376)
g32852(1) = NOT(g30614)
g34543(1) = NOT(g34359)
g32963(1) = NOT(g30825)
g32664(1) = NOT(g31528)
g32576(1) = NOT(g30614)
g32484(1) = NOT(g31566)
g32554(1) = NOT(g30614)
g32609(1) = NOT(g30735)
g32608(1) = NOT(g31376)
g32921(1) = NOT(g31672)
g32745(1) = NOT(g31376)
g32799(1) = NOT(g31710)
g32813(1) = NOT(g31710)
g32798(1) = NOT(g31672)
g32973(1) = NOT(g31021)
g32805(1) = NOT(g31672)
g32674(1) = NOT(g30735)
g32732(1) = NOT(g30825)
g32934(1) = NOT(g30735)
g32692(1) = NOT(g31528)
g32761(1) = NOT(g30825)
g32539(1) = NOT(g31170)
g32538(1) = NOT(g31070)
g32771(1) = NOT(g31021)
g32683(1) = NOT(g30614)
g32515(1) = NOT(g30825)
g32882(1) = NOT(g31376)
g32584(1) = NOT(g30673)
g32759(1) = NOT(g31376)
g32725(1) = NOT(g30825)
g32758(1) = NOT(g31327)
g32744(1) = NOT(g31327)
g32849(1) = NOT(g31021)
g32940(1) = NOT(g31376)
g32848(1) = NOT(g30825)
g32652(1) = NOT(g30735)
g32804(1) = NOT(g30735)
g32962(1) = NOT(g30735)
g32500(1) = NOT(g30735)
g32833(1) = NOT(g30825)
g34346(1) = NOT(g34162)
g32613(1) = NOT(g30673)
g32947(1) = NOT(g31376)
g32605(1) = NOT(g30614)
g32812(1) = NOT(g30825)
g32463(1) = NOT(g31566)
g32951(1) = NOT(g31021)
g32972(1) = NOT(g31710)
g32033(1) = NOT(g30929)
g32795(1) = NOT(g31327)
g32514(1) = NOT(g30735)
g32507(1) = NOT(g30735)
g32541(1) = NOT(g30673)
g32473(1) = NOT(g31070)
g32789(1) = NOT(g30735)
g32788(1) = NOT(g31327)
g32724(1) = NOT(g30735)
g32829(1) = NOT(g30937)
g32920(1) = NOT(g30825)
g32535(1) = NOT(g31554)
g32828(1) = NOT(g31710)
g32946(1) = NOT(g31327)
g32682(1) = NOT(g30825)
g32760(1) = NOT(g30735)
g32506(1) = NOT(g31376)
g32927(1) = NOT(g30825)
g32649(1) = NOT(g30673)
g32648(1) = NOT(g30614)
g32491(1) = NOT(g31566)
g32903(1) = NOT(g31376)
g32604(1) = NOT(g31154)
g32755(1) = NOT(g31672)
g32770(1) = NOT(g31710)
g32563(1) = NOT(g31554)
g32767(1) = NOT(g30735)
g32794(1) = NOT(g30937)
g32899(1) = NOT(g31021)
g32633(1) = NOT(g31154)
g32898(1) = NOT(g30825)
g32719(1) = NOT(g31672)
g32718(1) = NOT(g30825)
g32521(1) = NOT(g31376)
g32832(1) = NOT(g30735)
g32861(1) = NOT(g31376)
g32573(1) = NOT(g30825)
g32926(1) = NOT(g31376)
g32612(1) = NOT(g30614)
g32099(3) = NOT(g31009)
g32701(1) = NOT(g31376)
g32777(1) = NOT(g31710)
g32534(1) = NOT(g30673)
g32462(1) = NOT(g30673)
g32766(1) = NOT(g31376)
g32871(1) = NOT(g30937)
g32629(1) = NOT(g31376)
g30105(1) = NOT(I28336)
g32472(1) = NOT(g30825)
g32628(1) = NOT(g31542)
g32911(1) = NOT(g31376)
g32591(1) = NOT(g30614)
g32776(1) = NOT(g31672)
g32785(1) = NOT(g31710)
g32754(1) = NOT(g30825)
g32859(1) = NOT(g30614)
g32825(1) = NOT(g30735)
g32950(1) = NOT(g31672)
g32858(1) = NOT(g31327)
g32844(1) = NOT(g30937)
g33261(1) = OR(g32111, g29525)
g33393(1) = OR(g32286, g29984)
g32203(1) = AND(g4249, g31327)
g32281(1) = AND(g31257, g20500)
g32301(1) = AND(g31276, g20547)
g31273(1) = AND(g30143, g27779)
g33106(1) = AND(g32408, g18990)
g32290(1) = AND(g31267, g20525)
g32376(1) = AND(g2689, g31710)
g32095(1) = AND(g7619, g30825)
g32239(1) = OR(g30595, g29350)
g34310(1) = AND(g14003, g34162)
g29908(1) = NOR(g6918, g28471)
g32089(1) = AND(g27261, g31021)
g32088(1) = AND(g27241, g31070)
g32338(1) = AND(g31466, g20668)
g32315(1) = AND(g31306, g23517)
g32250(1) = OR(g30598, g29351)
g32055(1) = AND(g10999, g30825)
g32070(1) = AND(g10967, g30825)
g33271(1) = OR(g32120, g29549)
g31324(1) = AND(g30171, g27937)
g32067(1) = AND(g4727, g30614)
g31272(1) = AND(g30117, g27742)
g32196(1) = AND(g27587, g31376)
g32018(1) = AND(g4146, g30937)
g30316(1) = AND(g29199, g7097, g6682)
g32402(1) = AND(g4888, g30990)
g33281(1) = OR(g32142, g29576)
g32256(1) = AND(g31249, g20382)
g30273(1) = NOR(g5990, g29036)
g32300(1) = AND(g31274, g20544)
g33268(1) = OR(g32116, g29538)
g33257(1) = OR(g32108, g29519)
g32314(1) = AND(g31304, g23516)
g32287(1) = AND(g2823, g30578)
g32307(1) = AND(g31291, g23500)
g32085(1) = AND(g27253, g31021)
g32054(1) = AND(g10890, g30735)
g32269(1) = AND(g31253, g20443)
g31281(1) = AND(g30106, g27742)
g31301(1) = AND(g30170, g27907)
g32180(1) = AND(g2791, g31638)
g29898(1) = NOR(g6895, g28458)
g32335(1) = AND(g6199, g31566)
g32278(1) = AND(g2811, g30572)
g30282(1) = NOR(g6336, g29073)
g32306(1) = AND(g31289, g23499)
g30672(1) = OR(g13737, g29752)
g28683(1) = AND(g27876, g20649)
g34048(1) = NAND(g33669, g10583, g7442)
g31297(1) = AND(g30144, g27837)
g33303(1) = OR(g32159, g29638)
g30597(1) = OR(g13564, g29693)
g32410(1) = AND(g4933, g30997)
g34309(1) = AND(g13947, g34147)
g30308(1) = AND(g29178, g7004, g5297)
g32084(1) = AND(g10948, g30825)
g33270(1) = OR(g32119, g29547)
g32321(1) = AND(g27613, g31376)
g32179(1) = AND(g31748, g27907)
g32178(1) = AND(g31747, g27886)
g31987(1) = AND(g31767, g22198)
g31943(1) = AND(g4717, g30614)
g33384(1) = OR(g32248, g29943)
g31296(1) = AND(g30119, g27779)
g31968(1) = AND(g31757, g22168)
g33265(1) = OR(g32113, g29530)
g33280(1) = OR(g32141, g29574)
g33277(1) = OR(g32129, g29568)
g32266(1) = OR(g30604, g29354)
g32242(1) = AND(g31245, g20324)
g31496(1) = AND(g2338, g30312)
g31986(1) = AND(g31766, g22197)
g32293(1) = AND(g2827, g30593)
g32265(1) = AND(g2799, g30567)
g33287(1) = OR(g32146, g29586)
g29886(1) = NOR(g3288, g28458)
g32014(1) = AND(g8715, g30673)
g33276(1) = OR(g32128, g29566)
g32340(1) = AND(g31468, g23585)
g32035(1) = AND(g4176, g30937)
g29315(1) = AND(g29188, g7051, g5990)
g31300(1) = AND(g30148, g27858)
g34524(1) = AND(g9083, g34359)
g30290(1) = NOR(g6682, g29110)
g30732(1) = OR(g13778, g29762)
g33286(1) = OR(g32145, g29585)
g33296(1) = OR(g32156, g29617)
g32165(1) = AND(g31669, g27742)
g31480(1) = AND(g1644, g30296)
g31314(1) = AND(g30183, g27937)
g32175(1) = AND(g31709, g27858)
g31970(1) = NOR(g9024, g30583)
g33383(1) = OR(g32244, g29940)
I31593(1) = AND(g31003, g8350, g7788)
g29873(1) = NOR(g6875, g28458)
g31993(1) = AND(g31774, g22214)
I31600(1) = AND(g31009, g8400, g7809)
g31502(1) = AND(g2472, g29311)
g32274(1) = AND(g31256, g20447)
g31286(1) = AND(g30159, g27858)
g32292(1) = AND(g31269, g20530)
g31975(1) = AND(g31761, g22177)
g32409(1) = AND(g4754, g30996)
g28360(1) = AND(g27401, g19861)
g33295(1) = OR(g32153, g29605)
g30733(1) = OR(g13807, g29773)
g32283(1) = AND(g31259, g20506)
g32303(1) = AND(g27550, g31376)
g31321(1) = AND(g30146, g27886)
g32174(1) = AND(g31708, g27837)
g29900(1) = NOR(g3639, g28471)
g32225(1) = OR(g30576, g29336)
g32326(1) = AND(g31317, g23539)
g31242(1) = AND(g29373, g25409)
g32183(1) = AND(g2795, g31653)
g31974(1) = AND(g31760, g22176)
g33386(1) = OR(g32258, g29951)
g30285(1) = NOR(g7097, g29110)
g34330(1) = OR(g34069, g33717)
g31992(1) = AND(g31773, g22213)
g33254(1) = OR(g32104, g29512)
g32047(1) = AND(g27248, g31070)
g32311(1) = AND(g31295, g20582)
g31275(1) = AND(g30147, g27800)
g32350(1) = AND(g2697, g31710)
g31237(1) = AND(g29366, g25325)
g32396(1) = AND(g4698, g30983)
g32020(1) = AND(g4157, g30937)
g32046(1) = AND(g10925, g30735)
g33273(1) = OR(g32122, g29553)
g32282(1) = AND(g31258, g20503)
g32302(1) = AND(g31279, g23485)
g32105(1) = AND(g4922, g30673)
g31965(1) = NOR(g30583, g4358)
g30262(1) = NOR(g5644, g29008)
g32204(1) = AND(g4245, g31327)
g32356(1) = AND(g2704, g31710)
g32182(1) = AND(g31753, g27937)
g32331(1) = AND(g31322, g20637)
g29889(1) = NOR(g6905, g28471)
g34344(1) = AND(g34107, g20038)
g32097(1) = AND(g25960, g31021)
g32343(1) = AND(g31473, g20710)
g31283(1) = AND(g30156, g27837)
g32369(1) = AND(g2130, g31672)
g32412(1) = AND(g4765, g30998)
g29910(1) = NOR(g3990, g28484)
g33253(1) = OR(g32103, g29511)
g28660(1) = AND(g27824, g20623)
g32310(1) = AND(g27577, g31376)
g32050(1) = AND(g11003, g30825)
g33272(1) = OR(g32121, g29551)
g31949(1) = AND(g1287, g30825)
g30249(1) = NOR(g5297, g28982)
g33260(1) = OR(g32110, g29524)
g31933(1) = AND(g939, g30735)
g29903(1) = NOR(g6928, g28484)
g33282(1) = OR(g32143, g29577)
g32317(1) = AND(g5507, g31542)
g32323(1) = AND(g31311, g20610)
g31942(1) = NOR(g8977, g30583)
g32232(1) = AND(g31241, g20266)
g32261(1) = AND(g31251, g20386)
g33259(1) = OR(g32109, g29521)
g32056(1) = AND(g27271, g31021)
g32342(1) = AND(g6545, g31579)
g31282(1) = AND(g30130, g27779)
g30916(1) = OR(g13853, g29799)
g32198(1) = AND(g4253, g31327)
g33387(1) = OR(g32263, g29954)
g32330(1) = AND(g31320, g20631)
g33292(1) = OR(g32150, g29601)
g32161(1) = AND(g3151, g31154)
g32087(1) = AND(g1291, g30825)
g32069(1) = AND(g10878, g30735)
g28639(1) = AND(g27767, g20597)
g33390(1) = OR(g32276, g29968)
g32337(1) = AND(g31465, g20663)
g32171(1) = AND(g31706, g27800)
g30240(1) = NOR(g7004, g28982)
g31513(1) = AND(g2606, g29318)
g32010(1) = AND(g31785, g22303)
g31961(1) = AND(g31751, g22154)
g31505(1) = AND(g30195, g24379)
g32086(1) = AND(g7597, g30735)
g32322(1) = AND(g31308, g20605)
g32238(1) = OR(g30594, g29349)
g32295(1) = AND(g27931, g31376)
g33389(1) = OR(g32272, g29964)
g30288(1) = NOR(g7087, g29073)
g32309(1) = AND(g5160, g31528)
g32224(1) = AND(g4300, g31327)
g28703(1) = AND(g27925, g20680)
g31310(1) = AND(g30157, g27886)
g31959(1) = AND(g4907, g30673)
g31944(1) = AND(g31745, g22146)
g32260(1) = AND(g31250, g20385)
g30734(1) = OR(g13808, g29774)
g32231(1) = OR(g30590, g29346)
g33267(1) = OR(g32115, g29535)
g30315(1) = AND(g29182, g7028, g5644)
g32230(1) = OR(g30589, g29345)
g32042(1) = AND(g27244, g31070)
g32255(1) = AND(g31248, g20381)
g30824(1) = OR(g13833, g29789)
g32270(1) = AND(g31254, g20444)
g32188(1) = AND(g27586, g31376)
g31323(1) = AND(g30150, g27907)
g31299(1) = AND(g30123, g27800)
g32030(1) = AND(g4172, g30937)
g31298(1) = AND(g30169, g27886)
g30294(1) = NOR(g7110, g29110)
g33266(1) = OR(g32114, g29532)
g33290(1) = OR(g32149, g29589)
g28327(1) = AND(g27365, g19785)
g31989(1) = AND(g31770, g22200)
g31988(1) = AND(g31768, g22199)
g32419(1) = AND(g4955, g31000)
g32170(1) = AND(g31671, g27779)
g29323(1) = AND(g28539, g6905, g3639)
g33298(1) = OR(g32158, g29622)
g32167(1) = AND(g3853, g31194)
g33256(1) = OR(g32107, g29517)
g31960(1) = AND(g31749, g22153)
g33279(1) = OR(g32140, g29573)
g33278(1) = OR(g32139, g29572)
g32313(1) = AND(g31303, g23515)
g30276(1) = NOR(g7074, g29073)
g32305(1) = AND(g31287, g20567)
g29915(1) = NOR(g6941, g28484)
g29316(1) = AND(g28528, g6875, g3288)
g30608(1) = OR(g13604, g29736)
g33289(1) = OR(g32148, g29588)
g33288(1) = OR(g32147, g29587)
g33297(1) = OR(g32157, g29621)
g32009(1) = AND(g31782, g22224)
g31967(1) = AND(g31755, g22167)
g31994(1) = AND(g31775, g22215)
g32008(1) = AND(g31781, g22223)
g32176(1) = AND(g2779, g31623)
g31977(1) = AND(g31764, g22179)
g29539(1) = OR(g2864, g28220)
g31966(1) = AND(g31754, g22166)
g31309(1) = AND(g30132, g27837)
g32083(1) = AND(g947, g30735)
g32348(1) = AND(g2145, g31672)
g30280(1) = NOR(g7064, g29036)
g32284(1) = AND(g31260, g20507)
g32304(1) = AND(g31284, g20564)
g31495(1) = AND(g1913, g30309)
g31976(1) = AND(g31762, g22178)
g31985(1) = AND(g4722, g30614)
g29322(1) = AND(g29192, g7074, g6336)
g32333(1) = AND(g31326, g23559)
g33255(1) = OR(g32106, g29514)
g31489(1) = AND(g2204, g30305)
g31488(1) = AND(g1779, g30302)
g32312(1) = AND(g31302, g20591)
g32200(1) = AND(g27468, g31376)
g33275(1) = OR(g32127, g29564)
g30611(1) = OR(g13671, g29743)
g30265(1) = NOR(g7051, g29036)
g32400(1) = AND(g4743, g30989)
g32013(1) = AND(g8673, g30614)
g30271(1) = NOR(g7041, g29008)
g33251(1) = OR(g32096, g29509)
g32328(1) = AND(g5853, g31554)
g32241(1) = AND(g31244, g20323)
g31467(1) = AND(g30162, g27937)
g28343(1) = AND(g27380, g19799)
g34523(1) = AND(g9162, g34351)
g32414(1) = AND(g4944, g30999)
g31266(1) = AND(g30129, g27742)
g30609(1) = OR(g13633, g29742)
g32082(1) = AND(g4917, g30673)
g33274(1) = OR(g32126, g29563)
g31313(1) = AND(g30160, g27907)
g32345(1) = AND(g2138, g31672)
g31285(1) = AND(g30134, g27800)
g31935(1) = NOR(g30583, g4349)
g33101(1) = AND(g32398, g18976)
g32332(1) = AND(g31325, g23558)
g34542(1) = AND(g34332, g20089)
g32049(1) = AND(g10902, g30735)
g32273(1) = AND(g31255, g20446)
g31941(1) = AND(g1283, g30825)
g33380(1) = OR(g32234, g29926)
g33294(1) = OR(g32152, g29604)
g32163(1) = AND(g3502, g31170)
g31501(1) = AND(g2047, g29310)
g32325(1) = AND(g31316, g23538)
g28722(1) = AND(g27955, g20738)
g32427(1) = OR(g8928, g30583)
g32291(1) = AND(g31268, g20527)
g34537(1) = OR(g34324, g34084)
g31312(1) = AND(g30136, g27858)
g32191(1) = AND(g27593, g31376)
g30252(1) = NOR(g7028, g29008)
g32324(1) = AND(g31315, g23537)
g32098(1) = AND(g4732, g30614)
g31991(1) = AND(g4912, g30673)
g33293(1) = OR(g32151, g29602)
g32246(1) = AND(g31246, g20326)
g32251(1) = OR(g30599, g29352)
g30260(1) = NOR(g7018, g28982)
g32071(1) = AND(g27236, g31070)
g29328(1) = AND(g28553, g6928, g3990)
g32172(1) = AND(g2767, g31608)
g31940(1) = AND(g943, g30735)
g33262(1) = OR(g32112, g29528)
I30330(1) = OR(g29385, g31376, g30735, g30825)
g30613(1) = NOR(g4507, g29365)
g30317(1) = OR(g29208, I28566, I28567)
I30124(1) = OR(g31070, g31154, g30614, g30673)
I29986(1) = OR(g31070, g31194, g30614, g30673)
I28147(1) = OR(g2946, g24561, g28220)
I30400(1) = OR(g31021, g30937, g31327, g30614)
I30399(1) = OR(g29385, g31376, g30735, g30825)
I30262(1) = OR(g31672, g31710, g31021, g30937)
I30055(1) = OR(g31070, g31170, g30614, g30673)
I30054(1) = OR(g29385, g31376, g30735, g30825)
I30469(1) = OR(g31672, g31710, g31021, g30937)
I30468(1) = OR(g29385, g31376, g30735, g30825)
I30123(1) = OR(g29385, g31376, g30735, g30825)
I29985(1) = OR(g29385, g31376, g30735, g30825)
I30193(1) = OR(g31070, g30614, g30673, g31528)
I30192(1) = OR(g29385, g31376, g30735, g30825)
I30331(1) = OR(g31672, g31710, g31021, g30937)
I30261(1) = OR(g29385, g31376, g30735, g30825)
g31997(10) = NAND(g22306, g30580)
g29540(6) = NAND(g28336, g13464)
g31978(6) = NAND(g30580, g15591)
g29556(6) = NAND(g28349, g13486)
g31793(1) = OR(g28031, g30317)
g33064(1) = OR(g31993, g22067)
g33026(1) = OR(g32307, g21795)
g33022(1) = OR(g32306, g21750)
g33049(1) = OR(g31966, g21929)
g32997(1) = OR(g32269, g18378)
g33063(1) = OR(g31988, g22066)
g33541(1) = OR(g33101, g18223)
g29303(1) = OR(g28703, g18801)
g33013(1) = OR(g32283, g18484)
g32994(1) = OR(g32290, g18367)
g32996(1) = OR(g32256, g18377)
g33016(1) = OR(g32284, g18509)
g33029(1) = OR(g32332, g21798)
g33027(1) = OR(g32314, g21796)
g33024(1) = OR(g32324, g21752)
g33053(1) = OR(g31967, g21974)
g33008(1) = OR(g32261, g18457)
g32990(1) = OR(g32281, g18341)
g33059(1) = OR(g31987, g22021)
g33007(1) = OR(g32331, g18455)
g33058(1) = OR(g31976, g22020)
g33006(1) = OR(g32291, g18447)
g33033(1) = OR(g32333, g21843)
g33032(1) = OR(g32326, g21842)
g33060(1) = OR(g31992, g22022)
g33023(1) = OR(g32313, g21751)
g32991(1) = OR(g32322, g18349)
g29268(1) = OR(g28343, g18625)
g33017(1) = OR(g32292, g18510)
g33055(1) = OR(g31986, g21976)
g33018(1) = OR(g32312, g18525)
g33067(1) = OR(g31989, g22111)
g33034(1) = OR(g32340, g21844)
g33050(1) = OR(g31974, g21930)
g33015(1) = OR(g32343, g18507)
g31896(1) = OR(g31242, g24305)
g29309(1) = OR(g28722, g18818)
g33062(1) = OR(g31977, g22065)
g33009(1) = OR(g32273, g18458)
g32995(1) = OR(g32330, g18375)
g33057(1) = OR(g31968, g22019)
g33031(1) = OR(g32315, g21841)
g34439(1) = OR(g34344, g18181)
g33012(1) = OR(g32274, g18483)
g32989(1) = OR(g32241, g18326)
g33021(1) = OR(g32302, g21749)
g34599(1) = OR(g34542, g18149)
g29285(1) = OR(g28639, g18750)
g29262(1) = OR(g28327, g18608)
g33004(1) = OR(g32246, g18431)
g33054(1) = OR(g31975, g21975)
g33065(1) = OR(g32008, g22068)
g29291(1) = OR(g28660, g18767)
g33052(1) = OR(g31961, g21973)
g33003(1) = OR(g32323, g18429)
g31897(1) = OR(g31237, g24322)
g33014(1) = OR(g32305, g18499)
g32992(1) = OR(g32242, g18351)
g32998(1) = OR(g32300, g18393)
g32987(1) = OR(g32311, g18323)
g33070(1) = OR(g32010, g22114)
g32999(1) = OR(g32337, g18401)
g33005(1) = OR(g32260, g18432)
g33002(1) = OR(g32304, g18419)
g33048(1) = OR(g31960, g21928)
g29297(1) = OR(g28683, g18784)
g33069(1) = OR(g32009, g22113)
g29274(1) = OR(g28360, g18642)
g33000(1) = OR(g32270, g18403)
g31895(1) = OR(g31505, g24296)
g33068(1) = OR(g31994, g22112)
g33001(1) = OR(g32282, g18404)
g33047(1) = OR(g31944, g21927)
g33011(1) = OR(g32338, g18481)
g33010(1) = OR(g32301, g18473)
g32988(1) = OR(g32232, g18325)
g32993(1) = OR(g32255, g18352)
g33028(1) = OR(g32325, g21797)
g33543(1) = OR(g33106, g18281)
g32394(1) = NOT(g30601)
g32318(2) = NOT(g31596)
g32446(2) = NOT(g31596)
g32377(2) = NOT(g30984)
I27579(1) = NOT(g28184)
g32407(1) = NOT(I29939)
g29371(1) = NOT(I27735)
I27564(1) = NOT(g28166)
g32024(2) = NOT(I29582)
g29358(1) = NOT(I27718)
g31794(1) = NOT(I29368)
g34545(3) = NAND(g11679, g794, g34354)
g29491(2) = NOT(I27777)
I27552(1) = NOT(g28162)
I29894(1) = NOT(g31771)
I27576(1) = NOT(g28173)
g30295(1) = NOT(I28540)
g33127(1) = NOT(g31950)
g33385(1) = NOT(g32038)
g33354(1) = NOT(g32329)
I27742(1) = NOT(g28819)
I27549(1) = NOT(g28161)
I29965(1) = NOT(g31189)
g32442(2) = NOT(g31213)
I28390(1) = NOT(g29185)
g32430(2) = NOT(g30984)
I29909(1) = NOT(g31791)
I27561(1) = NOT(g28163)
g32021(2) = NOT(I29579)
g31487(1) = NOT(I29149)
I28883(1) = NOT(g30105)
g31479(1) = NOT(I29139)
g29498(2) = NOT(I27784)
I27546(1) = NOT(g29041)
I27558(1) = NOT(g28155)
I28866(1) = NOT(g29730)
I29913(1) = NOT(g30605)
I27567(1) = NOT(g28181)
g34539(1) = NOT(g34354)
I29199(1) = NOT(g30237)
I28838(1) = NOT(g29372)
I28925(1) = NOT(g29987)
g32421(2) = NOT(g31213)
g33142(1) = NOT(g32072)
I27555(1) = NOT(g28142)
I27570(1) = NOT(g28262)
I28908(1) = NOT(g30182)
I29977(1) = NOT(g31596)
g33136(1) = NOT(g32057)
I29961(1) = NOT(g30984)
g31945(2) = NOT(g31189)
g33413(1) = NOT(g31971)
I29973(1) = NOT(g31213)
g32393(1) = NOT(g30922)
g34169(1) = AND(g33804, g31227)
g34698(1) = NOT(g34550)
g30072(1) = NOT(I28301)
I27573(1) = NOT(g28157)
g29368(1) = NOT(I27730)
g29379(1) = NOT(I27749)
g30116(1) = NOT(I28349)
g29353(1) = NOT(I27713)
g33382(1) = NOT(g32033)
g32434(2) = NOT(g31189)
g33848(1) = AND(g33261, g20384)
g33652(1) = AND(g33393, g18889)
I31246(1) = AND(g31672, g31839, g32810, g32811)
g31127(1) = NOR(g4966, g29556)
I31071(1) = AND(g31170, g31808, g32557, g32558)
g32355(1) = OR(g29855, g31286)
I31147(1) = AND(g32668, g32669, g32670, g32671)
I31196(1) = AND(g30825, g31830, g32738, g32739)
I31197(1) = AND(g32740, g32741, g32742, g32743)
g33093(1) = NOR(g31997, g4601)
g31483(1) = NOR(g4899, g29725)
I31151(1) = AND(g30825, g31822, g32673, g32674)
I31172(1) = AND(g32703, g32704, g32705, g32706)
g34513(1) = AND(g9003, g34346)
I31011(1) = AND(g30735, g31797, g32471, g32472)
I31012(1) = AND(g32473, g32474, g32475, g32476)
I31227(1) = AND(g32784, g32785, g32786, g32787)
g33138(1) = NOR(g32287, g31514)
g31117(1) = NOR(g4991, g29556)
I31266(1) = AND(g31327, g31843, g32838, g32839)
I31267(1) = AND(g32840, g32841, g32842, g32843)
I31281(1) = AND(g30735, g31845, g32861, g32862)
I31231(1) = AND(g31376, g31836, g32789, g32790)
I31232(1) = AND(g32791, g32792, g32793, g32794)
I31301(1) = AND(g31327, g31849, g32889, g32890)
g32374(1) = OR(g29895, g31323)
I31146(1) = AND(g30735, g31821, g32666, g32667)
I31061(1) = AND(g30825, g31806, g32543, g32544)
I31062(1) = AND(g32545, g32546, g32547, g32548)
g33434(1) = AND(g32239, g29702)
g33090(1) = NOR(g31997, g4593)
I31226(1) = AND(g29385, g32781, g32782, g32783)
I31127(1) = AND(g32638, g32639, g32640, g32641)
g30925(1) = AND(g29908, g23309)
g33143(1) = NOR(g32293, g31518)
I31297(1) = AND(g32884, g32885, g32886, g32887)
I31181(1) = AND(g29385, g32716, g32717, g32718)
g33094(1) = NOR(g31950, g4639)
g31240(1) = AND(g14793, g30206)
I31152(1) = AND(g32675, g32676, g32677, g32678)
g33447(1) = NOR(g31978, g7643)
I31211(1) = AND(g31021, g31833, g32759, g32760)
g31119(1) = NOR(g7898, g29556)
I31126(1) = AND(g30673, g31818, g32636, g32637)
g33419(1) = NOR(g31978, g7627)
g33141(1) = NOR(g32099, g8400)
g33147(1) = NOR(g32090, g7788)
I31302(1) = AND(g32891, g32892, g32893, g32894)
I31296(1) = AND(g30937, g31848, g32882, g32883)
g33088(1) = NOR(g31997, g7224)
g33440(1) = AND(g32250, g29719)
g33861(1) = AND(g33271, g20502)
g33162(1) = NOR(g4859, g32072)
I31006(1) = AND(g31376, g31796, g32464, g32465)
I31007(1) = AND(g32466, g32467, g32468, g32469)
I31202(1) = AND(g32747, g32748, g32749, g32750)
I31257(1) = AND(g32826, g32827, g32828, g32829)
I31111(1) = AND(g31070, g31815, g32615, g32616)
g33871(1) = AND(g33281, g20546)
I31067(1) = AND(g32552, g32553, g32554, g32555)
g31220(1) = AND(g30273, g25202)
I31056(1) = AND(g30735, g31805, g32536, g32537)
I31057(1) = AND(g32538, g32539, g32540, g32541)
g33137(1) = NOR(g4849, g32072)
g33100(1) = NOR(g32172, g31188)
g33859(1) = AND(g33426, g10531)
g33858(1) = AND(g33268, g20448)
I31001(1) = AND(g29385, g32456, g32457, g32458)
I31077(1) = AND(g32566, g32567, g32568, g32569)
g33844(1) = AND(g33257, g20327)
I31256(1) = AND(g31021, g31841, g32824, g32825)
g32373(1) = OR(g29894, g31321)
I31102(1) = AND(g32603, g32604, g32605, g32606)
I31157(1) = AND(g32682, g32683, g32684, g32685)
g32385(1) = OR(g31480, g29938)
g34695(1) = OR(g34523, g34322)
I31066(1) = AND(g31070, g31807, g32550, g32551)
g33085(1) = NOR(g31978, g4311)
g30919(1) = AND(g29898, g23286)
I31287(1) = AND(g32870, g32871, g32872, g32873)
I31307(1) = AND(g32898, g32899, g32900, g32901)
I31076(1) = AND(g30614, g31809, g32564, g32565)
g32352(1) = OR(g29852, g31282)
I31341(1) = AND(g31710, g31856, g32947, g32948)
I31156(1) = AND(g31070, g31823, g32680, g32681)
g31226(1) = AND(g30282, g25218)
g31476(1) = NOR(g4709, g29697)
g33135(1) = NOR(g32090, g8350)
I31101(1) = AND(g30735, g31813, g32601, g32602)
g32187(1) = AND(g30672, g25287)
I31131(1) = AND(g31542, g31819, g32643, g32644)
g34364(1) = AND(g34048, g24366)
g33107(1) = NOR(g32180, g31223)
g33889(1) = AND(g33303, g20641)
g32168(1) = AND(g30597, g25185)
I31286(1) = AND(g30825, g31846, g32868, g32869)
I31306(1) = AND(g30614, g31850, g32896, g32897)
I31187(1) = AND(g32726, g32727, g32728, g32729)
g34687(1) = AND(g14181, g34543)
g33860(1) = AND(g33270, g20501)
I31182(1) = AND(g32719, g32720, g32721, g32722)
g33148(1) = NOR(g4854, g32072)
I31217(1) = AND(g32768, g32769, g32770, g32771)
g33943(1) = AND(g33384, g21609)
g31969(1) = AND(g31189, g22139)
g33855(1) = AND(g33265, g20441)
g33870(1) = AND(g33280, g20545)
g32361(1) = OR(g29869, g31300)
I31331(1) = AND(g30825, g31854, g32933, g32934)
I31332(1) = AND(g32935, g32936, g32937, g32938)
I31321(1) = AND(g31376, g31852, g32919, g32920)
I31186(1) = AND(g31376, g31828, g32724, g32725)
I31212(1) = AND(g32761, g32762, g32763, g32764)
g33867(1) = AND(g33277, g20529)
g33450(1) = AND(g32266, g29737)
g33174(1) = NOR(g8714, g32072)
g33134(1) = NOR(g7686, g32057)
I31176(1) = AND(g31579, g31827, g32708, g32709)
I31177(1) = AND(g32710, g32711, g32712, g32713)
I31216(1) = AND(g30937, g31834, g32766, g32767)
I31117(1) = AND(g32624, g32625, g32626, g32627)
g33437(1) = NOR(g31997, g10275)
g33877(1) = AND(g33287, g20563)
g30915(1) = AND(g29886, g24778)
I31242(1) = AND(g32805, g32806, g32807, g32808)
I31326(1) = AND(g30735, g31853, g32926, g32927)
I31327(1) = AND(g32928, g32929, g32930, g32931)
g32351(1) = OR(g29851, g31281)
g33866(1) = AND(g33276, g20528)
g33144(1) = NOR(g4664, g32057)
g31231(1) = AND(g30290, g25239)
g32193(1) = AND(g30732, g25410)
I31116(1) = AND(g31154, g31816, g32622, g32623)
g33876(1) = AND(g33286, g20562)
g33885(1) = AND(g33296, g20609)
I31041(1) = AND(g31566, g31803, g32513, g32514)
I31251(1) = AND(g31710, g31840, g32817, g32818)
I31252(1) = AND(g32819, g32820, g32821, g32822)
I31237(1) = AND(g32798, g32799, g32800, g32801)
I31142(1) = AND(g32661, g32662, g32663, g32664)
I31096(1) = AND(g31376, g31812, g32594, g32595)
I31097(1) = AND(g32596, g32597, g32598, g32599)
g33163(1) = NOR(g32099, g7809)
g33269(1) = AND(g31970, g15582)
g33942(1) = AND(g33383, g21608)
I31222(1) = AND(g32775, g32776, g32777, g32778)
g30914(1) = AND(g29873, g20887)
I31347(1) = AND(g32956, g32957, g32958, g32959)
I31132(1) = AND(g32645, g32646, g32647, g32648)
I31236(1) = AND(g30735, g31837, g32796, g32797)
I31206(1) = AND(g31710, g31832, g32752, g32753)
I31207(1) = AND(g32754, g32755, g32756, g32757)
I31351(1) = AND(g30937, g31858, g32961, g32962)
I31137(1) = AND(g32654, g32655, g32656, g32657)
I31042(1) = AND(g32515, g32516, g32517, g32518)
I31036(1) = AND(g30673, g31802, g32506, g32507)
I31037(1) = AND(g32508, g32509, g32510, g32511)
g33449(1) = NOR(g10311, g31950)
I31021(1) = AND(g31070, g31799, g32485, g32486)
g33884(1) = AND(g33295, g20590)
g32164(1) = AND(g30733, g25171)
g32360(1) = OR(g29868, g31299)
I31091(1) = AND(g29385, g32586, g32587, g32588)
I31092(1) = AND(g32589, g32590, g32591, g32592)
I31346(1) = AND(g31021, g31857, g32954, g32955)
I31122(1) = AND(g32631, g32632, g32633, g32634)
I31086(1) = AND(g31554, g31811, g32578, g32579)
I31087(1) = AND(g32580, g32581, g32582, g32583)
I31292(1) = AND(g32877, g32878, g32879, g32880)
I31136(1) = AND(g29385, g32651, g32652, g32653)
g33448(1) = NOR(g7785, g31950)
I31352(1) = AND(g32963, g32964, g32965, g32966)
g33125(1) = NOR(g8606, g32057)
g31936(1) = AND(g31213, g24005)
g32371(1) = OR(g29883, g31313)
g30921(1) = AND(g29900, g24789)
g33423(1) = AND(g32225, g29657)
g33131(1) = NOR(g4659, g32057)
g33092(1) = NOR(g31978, g4332)
I31192(1) = AND(g32733, g32734, g32735, g32736)
g33098(1) = NOR(g31997, g4616)
g31068(1) = NOR(g4801, g29540)
g33639(1) = AND(g33386, g18829)
g31230(1) = AND(g30285, g20751)
g32370(1) = OR(g29882, g31312)
g34538(1) = AND(g34330, g20054)
g33841(1) = AND(g33254, g20268)
I31247(1) = AND(g32812, g32813, g32814, g32815)
g32205(1) = AND(g30922, g28463)
g31506(1) = NOR(g4793, g29540)
g33161(1) = NOR(g32090, g7806)
I31161(1) = AND(g30614, g31824, g32687, g32688)
I31162(1) = AND(g32689, g32690, g32691, g32692)
I31022(1) = AND(g32487, g32488, g32489, g32490)
g33139(1) = NOR(g8650, g32057)
g31121(1) = NOR(g4776, g29540)
I31047(1) = AND(g32524, g32525, g32526, g32527)
I31282(1) = AND(g32863, g32864, g32865, g32866)
I31311(1) = AND(g30673, g31851, g32903, g32904)
I31051(1) = AND(g31376, g31804, g32529, g32530)
I31072(1) = AND(g32559, g32560, g32561, g32562)
I31312(1) = AND(g32905, g32906, g32907, g32908)
g33863(1) = AND(g33273, g20505)
I31046(1) = AND(g29385, g32521, g32522, g32523)
g33264(1) = AND(g31965, g21306)
g33108(1) = NOR(g32183, g31228)
I31276(1) = AND(g31376, g31844, g32854, g32855)
I31277(1) = AND(g32856, g32857, g32858, g32859)
I31357(1) = AND(g32970, g32971, g32972, g32973)
g32375(1) = OR(g29896, g31324)
g33095(1) = NOR(g31997, g7236)
g31208(1) = AND(g30262, g25188)
g33089(1) = NOR(g31978, g4322)
g32386(1) = OR(g31488, g29949)
I31027(1) = AND(g32494, g32495, g32496, g32497)
I31016(1) = AND(g30825, g31798, g32478, g32479)
I31017(1) = AND(g32480, g32481, g32482, g32483)
g32359(1) = OR(g29867, g31298)
g32358(1) = OR(g29866, g31297)
I31081(1) = AND(g30673, g31810, g32571, g32572)
g30920(1) = AND(g29889, g21024)
I31356(1) = AND(g31327, g31859, g32968, g32969)
g34506(1) = AND(g8833, g34354)
I31026(1) = AND(g31194, g31800, g32492, g32493)
g32392(1) = OR(g31513, g30000)
g30927(1) = AND(g29910, g24795)
g33840(1) = AND(g33253, g20267)
I31112(1) = AND(g32617, g32618, g32619, g32620)
g33862(1) = AND(g33272, g20504)
g33321(1) = OR(g29712, g32182)
g31133(1) = NOR(g7953, g29556)
g31183(1) = AND(g30249, g25174)
g33847(1) = AND(g33260, g20383)
I31241(1) = AND(g30825, g31838, g32803, g32804)
g30926(1) = AND(g29903, g21163)
g33872(1) = AND(g33282, g20548)
g33311(1) = AND(g31942, g12925)
I31317(1) = AND(g32914, g32915, g32916, g32917)
g33075(1) = NOR(g31997, g7163)
I31002(1) = AND(g32459, g32460, g32461, g32462)
g33846(1) = AND(g33259, g20380)
g32354(1) = OR(g29854, g31285)
I31261(1) = AND(g30937, g31842, g32831, g32832)
g33103(1) = NOR(g32176, g31212)
g31372(1) = NOR(g8796, g29697)
g32199(1) = AND(g30916, g25506)
g33640(1) = AND(g33387, g18831)
I31316(1) = AND(g29385, g32911, g32912, g32913)
g33881(1) = AND(g33292, g20586)
I31271(1) = AND(g29385, g32846, g32847, g32848)
I31342(1) = AND(g32949, g32950, g32951, g32952)
g33310(1) = OR(g29631, g32165)
I31031(1) = AND(g30614, g31801, g32499, g32500)
g31482(1) = NOR(g8883, g29697)
I31106(1) = AND(g30825, g31814, g32608, g32609)
I31107(1) = AND(g32610, g32611, g32612, g32613)
g31515(1) = NOR(g4983, g29556)
g32388(1) = OR(g31495, g29962)
g33130(1) = NOR(g32265, g31497)
g33647(1) = AND(g33390, g18878)
g31182(1) = AND(g30240, g20682)
I31262(1) = AND(g32833, g32834, g32835, g32836)
g33315(1) = OR(g29665, g32175)
I31221(1) = AND(g31327, g31835, g32773, g32774)
g32353(1) = OR(g29853, g31283)
I31337(1) = AND(g32942, g32943, g32944, g32945)
I31171(1) = AND(g31528, g31826, g32701, g32702)
g33433(1) = AND(g32238, g29694)
g33439(1) = NOR(g31950, g4633)
g33646(1) = AND(g33389, g18876)
g32336(1) = AND(g31596, g11842)
g32362(1) = OR(g29870, g31301)
I31322(1) = AND(g32921, g32922, g32923, g32924)
g34535(1) = OR(g34309, g34073)
g31229(1) = AND(g30288, g23949)
g33314(1) = OR(g29663, g32174)
I31336(1) = AND(g31672, g31855, g32940, g32941)
g33129(1) = NOR(g8630, g32072)
g32195(1) = AND(g30734, g25451)
g33097(1) = NOR(g31950, g4628)
g33429(1) = AND(g32231, g29676)
g33857(1) = AND(g33267, g20445)
g33428(1) = AND(g32230, g29672)
g33146(1) = NOR(g4669, g32057)
g32189(1) = AND(g30824, g25369)
g31232(1) = AND(g30294, g23972)
g33160(1) = NOR(g8672, g32057)
g33856(1) = AND(g33266, g20442)
g31261(1) = AND(g14754, g30259)
g33880(1) = AND(g33290, g20568)
I31191(1) = AND(g30735, g31829, g32731, g32732)
g33175(1) = NOR(g32099, g7828)
g31126(1) = NOR(g7928, g29540)
g33887(1) = AND(g33298, g20615)
g32194(1) = AND(g30601, g28436)
I31201(1) = AND(g31672, g31831, g32745, g32746)
g33843(1) = AND(g33256, g20325)
g31116(1) = NOR(g7892, g29540)
g33869(1) = AND(g33279, g20543)
g33868(1) = AND(g33278, g20542)
g31225(1) = AND(g30276, g21012)
I31052(1) = AND(g32531, g32532, g32533, g32534)
g32391(1) = OR(g31502, g29982)
g30930(1) = AND(g29915, g23342)
g31469(1) = NOR(g8822, g29725)
g32177(1) = AND(g30608, g25214)
I31167(1) = AND(g32696, g32697, g32698, g32699)
g33427(1) = NOR(g10278, g31950)
g33879(1) = AND(g33289, g20566)
g33878(1) = AND(g33288, g20565)
g33886(1) = AND(g33297, g20614)
g32380(1) = OR(g29907, g31467)
g33438(1) = NOR(g31950, g4621)
g32390(1) = OR(g31501, g29979)
I31166(1) = AND(g30673, g31825, g32694, g32695)
g33317(1) = OR(g29688, g32179)
g33128(1) = NOR(g4653, g32057)
g34685(1) = AND(g14164, g34550)
g31224(1) = AND(g30280, g23932)
g33132(1) = NOR(g4843, g32072)
g33842(1) = AND(g33255, g20322)
g32344(1) = OR(g29804, g31266)
I31141(1) = AND(g31376, g31820, g32659, g32660)
g33313(1) = OR(g29649, g32171)
g33865(1) = AND(g33275, g20526)
g31507(1) = NOR(g9064, g29556)
g32184(1) = AND(g30611, g25249)
g31219(1) = AND(g30265, g20875)
g31218(1) = AND(g30271, g23909)
g33837(1) = AND(g33251, g20233)
g33140(1) = NOR(g7693, g32072)
I31032(1) = AND(g32501, g32502, g32503, g32504)
g32372(1) = OR(g29884, g31314)
g33096(1) = NOR(g31997, g4608)
g32206(1) = AND(g30609, g25524)
g32349(1) = OR(g29840, g31275)
I31082(1) = AND(g32573, g32574, g32575, g32576)
g33864(1) = AND(g33274, g20524)
g33305(1) = AND(g31935, g17811)
g33432(1) = NOR(g31997, g6978)
g33316(1) = OR(g29685, g32178)
g33109(1) = NOR(g31997, g4584)
g33145(1) = NOR(g8677, g32072)
g31498(1) = NOR(g9030, g29540)
g33312(1) = OR(g29646, g32170)
I31121(1) = AND(g30614, g31817, g32629, g32630)
g32387(1) = OR(g31489, g29952)
g33941(1) = AND(g33380, g21560)
I31291(1) = AND(g31021, g31847, g32875, g32876)
g33883(1) = AND(g33294, g20589)
g33084(1) = NOR(g31978, g7655)
g33304(1) = AND(g32427, g31971)
g31318(1) = NOR(g4785, g29697)
g32368(1) = OR(g29881, g31310)
g34702(1) = AND(g34537, g20208)
g32347(1) = OR(g29839, g31273)
g31491(1) = NOR(g8938, g29725)
g31207(1) = AND(g30252, g20739)
g31373(1) = NOR(g4975, g29725)
I31272(1) = AND(g32849, g32850, g32851, g32852)
g33882(1) = AND(g33293, g20587)
g32367(1) = OR(g29880, g31309)
g32357(1) = OR(g29865, g31296)
g33441(1) = AND(g32251, g29722)
g31206(1) = AND(g30260, g23890)
g33133(1) = NOR(g32278, g31503)
g32389(1) = OR(g31496, g29966)
g33849(1) = AND(g33262, g20387)
g32346(1) = OR(g29838, g31272)
g32455(1) = NOR(g31566, I29985, I29986)
g32426(1) = OR(g26105, g26131, g30613)
I30728(1) = OR(g32345, g32350, g32056, g32018)
I30745(1) = OR(g31777, g32321, g32069, g32084)
I30746(1) = OR(g32047, g31985, g31991, g32309)
I30761(1) = OR(g32071, g32167, g32067, g32082)
g32845(1) = NOR(g30673, I30399, I30400)
g32780(1) = NOR(g31327, I30330, I30331)
I30740(1) = OR(g31776, g32188, g32083, g32087)
I30741(1) = OR(g32085, g32030, g32224, g32013)
I29351(1) = OR(g29328, g29323, g29316, g30316)
I30760(1) = OR(g31778, g32295, g32046, g32050)
I30755(1) = OR(g30564, g32303, g32049, g32055)
I30718(1) = OR(g32348, g32356, g32097, g32020)
g32585(1) = NOR(g31542, I30123, I30124)
g32520(1) = NOR(g31554, I30054, I30055)
I30727(1) = OR(g31759, g32196, g31933, g31941)
g32910(1) = NOR(g31327, I30468, I30469)
I30735(1) = OR(g32369, g32376, g32089, g32035)
I30750(1) = OR(g31788, g32310, g32054, g32070)
I30751(1) = OR(g32042, g32161, g31943, g31959)
I30734(1) = OR(g31790, g32191, g32086, g32095)
I30756(1) = OR(g32088, g32163, g32098, g32105)
I30717(1) = OR(g31787, g32200, g31940, g31949)
I29352(1) = OR(g29322, g29315, g30315, g30308)
g29914(1) = OR(g22531, g22585, I28147)
g32715(1) = NOR(g31327, I30261, I30262)
g32650(1) = NOR(g31579, I30192, I30193)
g33083(1) = NAND(g7805, g32118)
g29210(1) = NOT(I27546)
g29211(1) = NOT(I27549)
g29212(1) = NOT(I27552)
g29213(1) = NOT(I27555)
g29214(1) = NOT(I27558)
g29215(1) = NOT(I27561)
g29216(1) = NOT(I27564)
g29217(1) = NOT(I27567)
g29218(1) = NOT(I27570)
g29219(1) = NOT(I27573)
g29220(1) = NOT(I27576)
g29221(1) = NOT(I27579)
g32429(1) = OR(g30318, g31794)
g33982(1) = OR(g33865, g18372)
g34007(1) = OR(g33640, g18467)
g33974(1) = OR(g33846, g18345)
g33966(1) = OR(g33837, g18318)
g33973(1) = OR(g33840, g18344)
g33043(1) = OR(g32195, g24325)
g34015(1) = OR(g33858, g18502)
g34001(1) = OR(g33844, g18450)
g33976(1) = OR(g33869, g18347)
g33997(1) = OR(g33871, g18427)
g33042(1) = OR(g32193, g24324)
g33972(1) = OR(g33941, g18335)
g33993(1) = OR(g33646, g18413)
g33036(1) = OR(g32168, g24309)
g34014(1) = OR(g33647, g18493)
g33975(1) = OR(g33860, g18346)
g33037(1) = OR(g32177, g24310)
g33039(1) = OR(g32187, g24312)
g34003(1) = OR(g33866, g18452)
g33989(1) = OR(g33870, g18398)
g34005(1) = OR(g33883, g18454)
g33984(1) = OR(g33881, g18374)
g33967(1) = OR(g33842, g18319)
g34004(1) = OR(g33879, g18453)
g33990(1) = OR(g33882, g18399)
g34021(1) = OR(g33652, g18519)
g33969(1) = OR(g33864, g18321)
g34440(1) = OR(g34364, g24226)
g33038(1) = OR(g32184, g24311)
g34724(1) = OR(g34702, g18152)
g33991(1) = OR(g33885, g18400)
g33045(1) = OR(g32206, g24328)
g33970(1) = OR(g33868, g18322)
g34009(1) = OR(g33863, g18477)
g34018(1) = OR(g33887, g18505)
g34600(1) = OR(g34538, g18182)
g33988(1) = OR(g33861, g18397)
g34008(1) = OR(g33849, g18476)
g34012(1) = OR(g33886, g18480)
g34017(1) = OR(g33880, g18504)
g33983(1) = OR(g33877, g18373)
g33980(1) = OR(g33843, g18370)
g34011(1) = OR(g33884, g18479)
g33996(1) = OR(g33862, g18426)
g33995(1) = OR(g33848, g18425)
g34000(1) = OR(g33943, g18441)
g34016(1) = OR(g33867, g18503)
g33998(1) = OR(g33878, g18428)
g33977(1) = OR(g33876, g18348)
g34010(1) = OR(g33872, g18478)
g33986(1) = OR(g33639, g18387)
g33968(1) = OR(g33855, g18320)
g33994(1) = OR(g33841, g18424)
g34002(1) = OR(g33857, g18451)
g33979(1) = OR(g33942, g18361)
g33040(1) = OR(g32164, g24313)
g33041(1) = OR(g32189, g24323)
g33044(1) = OR(g32199, g24327)
g34019(1) = OR(g33889, g18506)
g33987(1) = OR(g33847, g18396)
g33981(1) = OR(g33856, g18371)
g33204(7) = OR(g32317, I30750, I30751)
I28594(1) = NOT(g29379)
g30729(1) = NOT(I28883)
I30901(1) = NOT(g32407)
g33187(9) = OR(g32014, I30740, I30741)
g33219(7) = OR(g32335, I30760, I30761)
g33197(6) = OR(g32342, I30745, I30746)
g31591(4) = OR(g29358, g29353)
g34697(1) = NOT(g34545)
g32381(1) = NOT(I29909)
g33164(9) = OR(g32203, I30727, I30728)
g32132(4) = OR(g31487, g31479)
I28591(1) = NOT(g29371)
g30991(4) = NOT(I28925)
g33176(9) = OR(g32198, I30734, I30735)
g33212(6) = OR(g32328, I30755, I30756)
I31791(1) = NOT(g33354)
I28872(1) = NOT(g30072)
g33149(9) = OR(g32204, I30717, I30718)
g30155(1) = NOT(I28390)
g30606(1) = NOT(I28866)
g32437(1) = NOT(I29965)
I29233(1) = NOT(g30295)
g33076(2) = OR(g32336, g32446)
I30962(1) = NOT(g32021)
I29248(1) = NOT(g29491)
I29236(1) = NOT(g29498)
g29374(1) = NOT(I27742)
I28588(1) = NOT(g29368)
g31578(1) = NOT(I29199)
g32383(1) = NOT(I29913)
g33430(1) = NOT(g32421)
I32352(1) = NOT(g34169)
g33323(2) = OR(g31936, g32442)
g32449(1) = NOT(I29977)
g32433(1) = NOT(I29961)
g33326(1) = NOT(g32318)
I30644(1) = NOT(g32024)
g34703(2) = NOR(g8899, g34545, g11083)
g33072(1) = NOT(g31945)
g32445(1) = NOT(I29973)
I29245(1) = NOT(g29491)
g32364(2) = NOT(I29894)
g30928(1) = NOT(I28908)
g31783(1) = OR(I29351, I29352)
I29239(1) = NOT(g29498)
I28582(1) = NOT(g30116)
g33375(1) = NOT(g32377)
g33318(2) = OR(g31969, g32434)
I30641(1) = NOT(g32024)
g30569(2) = NOT(I28838)
g33838(1) = NAND(g33083, g4369)
I30959(1) = NOT(g32021)
g33263(1) = AND(g32393, g25481)
g32420(1) = AND(g31127, g19533)
g33706(1) = OR(g32412, g33440)
g33406(1) = AND(g32355, g21399)
g33500(1) = AND(g32744, I31196, I31197)
g33833(1) = AND(g33093, g25852)
g32044(1) = AND(g31483, g20085)
g33463(1) = AND(g32477, I31011, I31012)
g32280(1) = OR(g24790, g31225)
g33795(1) = AND(g33138, g20782)
g32403(1) = AND(g31117, g15842)
g33514(1) = AND(g32844, I31266, I31267)
g33507(1) = AND(g32795, I31231, I31232)
g33421(1) = AND(g32374, g21455)
g33473(1) = AND(g32549, I31061, I31062)
g32252(1) = OR(g31183, g31206)
g33828(1) = AND(g33090, g24411)
g33760(1) = AND(g33143, g20328)
g33506(1) = AND(g32788, I31226, I31227)
g34742(1) = AND(g9000, g34698)
g33927(1) = AND(g33094, g21412)
g33491(1) = AND(g32679, I31151, I31152)
g33903(1) = AND(g33447, g19146)
g32411(1) = AND(g31119, g13469)
g33898(1) = AND(g33419, g15655)
g33719(1) = AND(g33141, g19433)
g33718(1) = AND(g33147, g19432)
g33521(1) = AND(g32895, I31301, I31302)
g33832(1) = AND(g33088, g27991)
g32130(1) = OR(g30921, g30925)
g33701(1) = AND(g33162, g16305)
g33462(1) = AND(g32470, I31006, I31007)
g31288(1) = OR(g2955, g29914)
g32253(1) = OR(g24771, g31207)
g33472(1) = AND(g32542, I31056, I31057)
g33911(1) = AND(g33137, g10725)
g33785(1) = AND(g33100, g20550)
g32279(1) = OR(g31220, g31224)
g33420(1) = AND(g32373, g21454)
g33446(1) = AND(g32385, g21607)
g34774(1) = AND(g34695, g20180)
g33902(1) = AND(g33085, g13202)
g33703(1) = OR(g32410, g33434)
g33699(1) = OR(g32409, g33433)
g32268(1) = OR(g24785, g31219)
g33403(1) = AND(g32352, g21396)
g32039(1) = AND(g31476, g20070)
g33715(1) = AND(g33135, g19416)
g33481(1) = AND(g32607, I31101, I31102)
g33490(1) = AND(g32672, I31146, I31147)
g33784(1) = AND(g33107, g20531)
g32294(1) = OR(g31231, g31232)
g33520(1) = AND(g32888, I31296, I31297)
g33497(1) = AND(g32723, I31181, I31182)
g34762(1) = OR(g34687, g34524)
g33700(1) = AND(g33148, g11012)
g33411(1) = AND(g32361, g21410)
g33527(1) = AND(g32939, I31331, I31332)
g34679(1) = AND(g14093, g34539)
g33503(1) = AND(g32765, I31211, I31212)
g33707(1) = AND(g33174, g13346)
g33910(1) = AND(g33134, g7836)
g33496(1) = AND(g32714, I31176, I31177)
g33111(1) = AND(g24005, g32421)
g33801(1) = AND(g33437, g25327)
g33692(1) = OR(g32400, g33428)
g33526(1) = AND(g32932, I31326, I31327)
g33402(1) = AND(g32351, g21395)
g33689(1) = AND(g33144, g11006)
g33511(1) = AND(g32823, I31251, I31252)
g33480(1) = AND(g32600, I31096, I31097)
g33721(1) = AND(g33163, g19440)
g32124(1) = OR(g24488, g30920)
g33734(1) = AND(g7806, g33136, I31593)
g33685(1) = OR(g32396, g33423)
g33487(1) = AND(g32649, I31131, I31132)
g33502(1) = AND(g32758, I31206, I31207)
g33469(1) = AND(g32519, I31041, I31042)
g33468(1) = AND(g32512, I31036, I31037)
g33815(1) = AND(g33449, g12911)
g33410(1) = AND(g32360, g21409)
g33714(1) = OR(g32419, g33450)
g33479(1) = AND(g32593, I31091, I31092)
g33478(1) = AND(g32584, I31086, I31087)
g33486(1) = AND(g32642, I31126, I31127)
g33922(1) = AND(g33448, g7202)
g33531(1) = AND(g32967, I31351, I31352)
g33676(1) = AND(g33125, g7970)
g32288(1) = OR(g31226, g31229)
g33417(1) = AND(g32371, g21424)
g33909(1) = AND(g33131, g10708)
g33908(1) = AND(g33092, g18935)
g32123(1) = OR(g30915, g30919)
g33814(1) = AND(g33098, g28144)
g32397(1) = AND(g31068, g15830)
g33112(1) = NOR(g31240, g32194)
g33416(1) = AND(g32370, g21423)
g33510(1) = AND(g32816, I31246, I31247)
g33835(1) = AND(g4340, g33413)
g34693(1) = OR(g34513, g34310)
g32051(1) = AND(g31506, g10831)
g33720(1) = AND(g33161, g19439)
g33493(1) = AND(g32693, I31161, I31162)
g33465(1) = AND(g32491, I31021, I31022)
g33237(1) = AND(g32394, g25198)
g33684(1) = AND(g33139, g13565)
g32413(1) = AND(g31121, g19518)
g33517(1) = AND(g32867, I31281, I31282)
g33709(1) = OR(g32414, g33441)
g33523(1) = AND(g32909, I31311, I31312)
g33475(1) = AND(g32563, I31071, I31072)
g33790(1) = AND(g33108, g20643)
g33516(1) = AND(g32860, I31276, I31277)
g33422(1) = AND(g32375, g21456)
g33834(1) = AND(g33095, g29172)
g33905(1) = AND(g33089, g15574)
g33073(1) = AND(g32386, g18828)
g33530(1) = AND(g32960, I31346, I31347)
g33464(1) = AND(g32484, I31016, I31017)
g33409(1) = AND(g32359, g21408)
g33408(1) = AND(g32358, g21407)
g33474(1) = AND(g32556, I31066, I31067)
g33492(1) = AND(g32686, I31156, I31157)
g33381(1) = AND(g11842, g32318)
g33091(1) = AND(g32392, g18897)
g33117(1) = NOR(g31261, g32205)
g33522(1) = AND(g32902, I31306, I31307)
g33483(1) = AND(g32621, I31111, I31112)
g33904(1) = AND(g33321, g21059)
g32428(1) = AND(g31133, g16261)
g33509(1) = AND(g32809, I31241, I31242)
g33508(1) = AND(g32802, I31236, I31237)
g33820(1) = AND(g33075, g26830)
g33405(1) = AND(g32354, g21398)
g34067(1) = NOR(g33859, g11772)
g33787(1) = AND(g33103, g20595)
g32031(1) = AND(g31372, g13464)
g33890(1) = AND(g33310, g20659)
g32144(1) = OR(g30927, g30930)
g32043(1) = AND(g31482, g16173)
g33482(1) = AND(g32614, I31106, I31107)
g32131(1) = OR(g24495, g30926)
g32068(1) = AND(g31515, g10862)
g33081(1) = AND(g32388, g18875)
g33786(1) = AND(g33130, g20572)
g33914(1) = OR(g33305, g33311)
g33513(1) = AND(g32837, I31261, I31262)
g33897(1) = AND(g33315, g20777)
g33505(1) = AND(g32779, I31221, I31222)
g33404(1) = AND(g32353, g21397)
g33811(1) = AND(g33439, g17573)
g33891(1) = OR(g33264, g33269)
g33412(1) = AND(g32362, g21411)
g34700(1) = AND(g34535, g20129)
g33896(1) = AND(g33314, g20771)
g33742(1) = AND(g7828, g33142, I31600)
g33681(1) = AND(g33129, g7991)
g33802(1) = AND(g33097, g14545)
g33730(1) = AND(g7202, g4621, g33127, g4633)
g33690(1) = AND(g33146, g16280)
g33504(1) = AND(g32772, I31216, I31217)
g33697(1) = AND(g33160, g13330)
g33512(1) = AND(g32830, I31256, I31257)
g33499(1) = AND(g32737, I31191, I31192)
g33498(1) = AND(g32730, I31186, I31187)
g33722(1) = AND(g33175, g19445)
g32418(1) = AND(g31126, g16239)
g33461(1) = AND(g32463, I31001, I31002)
g33529(1) = AND(g32953, I31341, I31342)
g33528(1) = AND(g32946, I31336, I31337)
g32401(1) = AND(g31116, g13432)
g33694(1) = OR(g32402, g33429)
g32267(1) = OR(g31208, g31218)
g33471(1) = AND(g32535, I31051, I31052)
g33087(1) = AND(g32391, g18888)
g32036(1) = AND(g31469, g13486)
g33810(1) = AND(g33427, g12768)
g33425(1) = AND(g32380, g21466)
g33919(1) = AND(g33438, g10795)
g33086(1) = AND(g32390, g18887)
g33532(1) = AND(g32974, I31356, I31357)
g33901(1) = AND(g33317, g20920)
g32240(1) = OR(g24757, g31182)
g33680(1) = AND(g33128, g4688)
g33495(1) = AND(g32707, I31171, I31172)
g33687(1) = AND(g33132, g4878)
g32289(1) = OR(g24796, g31230)
g33392(1) = AND(g32344, g21362)
g33489(1) = AND(g32665, I31141, I31142)
g33525(1) = AND(g32925, I31321, I31322)
g33488(1) = AND(g32658, I31136, I31137)
g33830(1) = AND(g33382, g20166)
g33893(1) = AND(g33313, g20706)
g32052(1) = AND(g31507, g13885)
g34684(1) = AND(g14178, g34545)
g33470(1) = AND(g32528, I31046, I31047)
g33915(1) = AND(g33140, g7846)
g33467(1) = AND(g32505, I31031, I31032)
g33494(1) = AND(g32700, I31166, I31167)
g33418(1) = AND(g32372, g21425)
g33822(1) = AND(g33385, g20157)
g33524(1) = AND(g32918, I31316, I31317)
g33836(1) = AND(g33096, g27020)
g33401(1) = AND(g32349, g21381)
g33477(1) = AND(g32577, I31081, I31082)
g33809(1) = AND(g33432, g30184)
g33900(1) = AND(g33316, g20913)
g33466(1) = AND(g32498, I31026, I31027)
g33808(1) = AND(g33109, g22161)
g33693(1) = AND(g33145, g13594)
g32048(1) = AND(g31498, g13869)
g33892(1) = AND(g33312, g20701)
g33476(1) = AND(g32570, I31076, I31077)
g33485(1) = AND(g32635, I31121, I31122)
g33074(1) = AND(g32387, g18830)
g32117(1) = OR(g24482, g30914)
g33519(1) = AND(g32881, I31291, I31292)
g33518(1) = AND(g32874, I31286, I31287)
g33501(1) = AND(g32751, I31201, I31202)
g33906(1) = AND(g33084, g22311)
g32029(1) = AND(g31318, g16482)
g33415(1) = AND(g32368, g21422)
g33484(1) = AND(g32628, I31116, I31117)
g33400(1) = AND(g32347, g21380)
g32045(1) = AND(g31491, g16187)
g32032(1) = AND(g31373, g16515)
g33515(1) = AND(g32853, I31271, I31272)
g33414(1) = AND(g32367, g21421)
g33407(1) = AND(g32357, g21406)
g33114(1) = AND(g22139, g31945)
g33758(1) = AND(g33133, g20269)
g33082(1) = AND(g32389, g18877)
g33399(1) = AND(g32346, g21379)
g33394(4) = NAND(g10159, g4474, g32426)
g30327(1) = NOT(I28582)
g30329(1) = NOT(I28588)
g30330(1) = NOT(I28591)
g30331(1) = NOT(I28594)
g31656(1) = NOT(I29236)
g31665(1) = NOT(I29245)
g33079(1) = NOT(I30641)
g33435(1) = NOT(I30959)
g33554(1) = OR(g33407, g18353)
g34036(1) = OR(g33722, g18715)
g34026(1) = OR(g33715, g18682)
g33560(1) = OR(g33404, g18369)
g34790(1) = OR(g34774, g18151)
g34034(1) = OR(g33719, g18713)
g33963(1) = OR(g33830, g18124)
g34035(1) = OR(g33721, g18714)
g33584(1) = OR(g33406, g18449)
g33593(1) = OR(g33417, g18482)
g33552(1) = OR(g33400, g18343)
g33971(1) = OR(g33890, g18330)
g34025(1) = OR(g33927, g18672)
g33962(1) = OR(g33822, g18123)
g33999(1) = OR(g33893, g18436)
g33601(1) = OR(g33422, g18508)
g33978(1) = OR(g33892, g18356)
g33985(1) = OR(g33896, g18382)
g33575(1) = OR(g33086, g18420)
g33553(1) = OR(g33403, g18350)
g33602(1) = OR(g33425, g18511)
g33559(1) = OR(g33073, g18368)
g33607(1) = OR(g33091, g18526)
g33562(1) = OR(g33414, g18379)
g34028(1) = OR(g33720, g18684)
g33546(1) = OR(g33402, g18327)
g33583(1) = OR(g33074, g18448)
g33569(1) = OR(g33415, g18402)
g34027(1) = OR(g33718, g18683)
g33600(1) = OR(g33418, g18501)
g33561(1) = OR(g33408, g18376)
g33576(1) = OR(g33401, g18423)
g34006(1) = OR(g33897, g18462)
g34020(1) = OR(g33904, g18514)
g33594(1) = OR(g33421, g18485)
g33591(1) = OR(g33082, g18474)
g34725(1) = OR(g34700, g18183)
g33570(1) = OR(g33420, g18405)
g33567(1) = OR(g33081, g18394)
g33585(1) = OR(g33411, g18456)
g33578(1) = OR(g33410, g18433)
g33544(1) = OR(g33392, g18317)
g33551(1) = OR(g33446, g18342)
g34013(1) = OR(g33901, g18488)
g33545(1) = OR(g33399, g18324)
g33577(1) = OR(g33405, g18430)
g33592(1) = OR(g33412, g18475)
g33586(1) = OR(g33416, g18459)
g33599(1) = OR(g33087, g18500)
g33616(1) = OR(g33237, g24314)
g33617(1) = OR(g33263, g24326)
g33992(1) = OR(g33900, g18408)
g33568(1) = OR(g33409, g18395)
I31776(1) = NOT(g33204)
I29447(1) = NOT(g30729)
I31786(1) = NOT(g33197)
I31515(1) = NOT(g33187)
I31482(1) = NOT(g33204)
I31610(1) = NOT(g33149)
I31497(1) = NOT(g33187)
I31694(1) = NOT(g33176)
I31659(1) = NOT(g33219)
I31625(1) = NOT(g33197)
g32450(2) = NOT(g31591)
I31796(1) = NOT(g33176)
g31666(1) = NOT(I29248)
I30686(1) = NOT(g32381)
I31581(1) = NOT(g33164)
I31619(1) = NOT(g33212)
g34345(1) = NOT(I32352)
g33451(2) = NOT(g32132)
I29969(1) = NOT(g30991)
g33831(1) = AND(g23088, g33149, g9104)
I31597(1) = NOT(g33187)
g33728(1) = AND(g22626, g10851, g33187)
g33377(1) = NOT(I30901)
I31550(1) = NOT(g33204)
I31539(1) = NOT(g33212)
g33346(2) = NOT(g32132)
I29891(1) = NOT(g31578)
I29571(1) = NOT(g31783)
I31807(1) = NOT(g33149)
g33080(1) = NOT(I30644)
I31486(1) = NOT(g33197)
g30610(1) = NOT(I28872)
g33674(1) = AND(g33164, g10710, g22319)
g33819(1) = AND(g23088, g33176, g9104)
I31800(1) = NOT(g33164)
I31569(1) = NOT(g33197)
g33695(1) = NOT(g33187)
I31814(1) = NOT(g33149)
I31779(1) = NOT(g33212)
g33923(1) = NOT(I31791)
I29936(1) = NOT(g30606)
I31523(1) = NOT(g33187)
I31586(1) = NOT(g33149)
g33683(1) = AND(g33149, g10727, g22332)
I30986(1) = NOT(g32437)
g31655(1) = NOT(I29233)
I31504(1) = NOT(g33164)
I31727(1) = NOT(g33076)
I30861(1) = NOT(g32383)
I31686(1) = NOT(g33164)
I29981(1) = NOT(g31591)
g31937(2) = NOT(g30991)
I31823(1) = NOT(g33149)
I31607(1) = NOT(g33164)
I28597(1) = NOT(g29374)
I31474(1) = NOT(g33212)
I31642(1) = NOT(g33204)
I31820(1) = NOT(g33323)
I31622(1) = NOT(g33204)
I31564(1) = NOT(g33204)
I31650(1) = NOT(g33212)
g33678(1) = AND(g33149, g10710, g22319)
I31803(1) = NOT(g33176)
g33436(1) = NOT(I30962)
I31672(1) = NOT(g33149)
I30980(1) = NOT(g32132)
I29444(1) = NOT(g30928)
g34208(1) = NOT(g33838)
I31545(1) = NOT(g33219)
I31770(1) = NOT(g33197)
g34766(1) = NOT(g34703)
I31528(1) = NOT(g33219)
g33675(1) = AND(g33164, g10727, g22332)
I31810(1) = NOT(g33164)
g33913(1) = AND(g23088, g33204, g9104)
I31459(1) = NOT(g33219)
I31817(1) = NOT(g33323)
I31701(1) = NOT(g33164)
I31561(1) = NOT(g33197)
g33704(1) = AND(g33176, g10710, g22319)
g33812(1) = AND(g23088, g33187, g9104)
g33725(1) = AND(g22626, g10851, g33176)
I28897(1) = NOT(g30155)
I30992(1) = NOT(g32445)
I30983(1) = NOT(g32433)
I31782(1) = NOT(g33219)
g33907(1) = AND(g23088, g33219, g9104)
I31555(1) = NOT(g33212)
g31657(1) = NOT(I29239)
I31616(1) = NOT(g33219)
I30995(1) = NOT(g32449)
I31466(1) = NOT(g33318)
g32438(2) = NOT(g30991)
g32415(2) = NOT(g31591)
g33686(1) = NOT(g33187)
I31724(1) = NOT(g33076)
I31500(1) = NOT(g33176)
I31463(1) = NOT(g33318)
g33921(1) = AND(g33187, g9104, g19200)
g33711(1) = AND(g33176, g10727, g22332)
I31604(1) = NOT(g33176)
g34081(1) = AND(g33706, g19552)
g34158(1) = OR(g33784, g19740)
g33371(1) = AND(g32280, g21155)
g33359(1) = AND(g32252, g20853)
g33240(1) = OR(g32052, g32068)
g33247(1) = AND(g32130, g19980)
g33360(1) = AND(g32253, g20869)
g34103(1) = OR(g33701, g33707)
g34189(1) = OR(g33801, g33808)
g34149(1) = OR(g33760, g19674)
g33370(1) = AND(g32279, g21139)
g34095(1) = OR(g33681, g33687)
g33925(1) = NAND(g33394, g4462, g4467)
g34079(1) = AND(g33703, g19532)
g34078(1) = AND(g33699, g19531)
g33366(1) = AND(g32268, g21010)
g34057(1) = OR(g33911, g33915)
g33376(1) = AND(g32294, g21268)
g34842(1) = AND(g34762, g20168)
g33236(1) = OR(g32044, g32045)
g33118(1) = OR(g32413, g32418)
g34075(1) = AND(g33692, g19517)
g34199(1) = OR(g33820, g33828)
g33243(1) = AND(g32124, g19947)
g33431(1) = AND(g32364, g32377)
g34074(1) = AND(g33685, g19498)
g34167(1) = OR(g33786, g19768)
g34083(1) = AND(g33714, g19573)
g34046(1) = OR(g33906, g33908)
g34207(1) = OR(g33835, g33304)
g33373(1) = AND(g32288, g21205)
g33242(1) = AND(g32123, g19931)
g33807(1) = AND(g33112, g25452)
g34771(1) = AND(g34693, g20147)
g34206(1) = OR(g33834, g33836)
g34082(1) = AND(g33709, g19554)
g33115(1) = OR(g32397, g32401)
g33238(1) = OR(g32048, g32051)
g34055(1) = OR(g33909, g33910)
g33679(1) = NAND(g33394, g10737, g10308)
g33796(1) = AND(g33117, g25267)
g34193(1) = OR(g33809, g33814)
g34170(1) = OR(g33790, g19855)
g33116(1) = OR(g32403, g32411)
g34370(1) = AND(g34067, g10554)
g34190(1) = OR(g33802, g33810)
g33119(1) = OR(g32420, g32428)
g33231(1) = OR(g32032, g32036)
g34043(1) = OR(g33903, g33905)
g34064(1) = OR(g33919, g33922)
g33930(1) = NAND(g33394, g12767, g9848)
g33249(1) = AND(g32144, g20026)
g33248(1) = AND(g32131, g19996)
g34226(1) = AND(g33914, g21467)
g34168(1) = OR(g33787, g19784)
g34211(1) = AND(g33891, g21349)
g34099(1) = OR(g33684, g33689)
g33379(1) = AND(g30984, g32364)
g34826(1) = OR(g34742, g34685)
g34741(1) = AND(g8899, g34697)
g31995(1) = AND(g28274, g30569)
g34066(1) = AND(g33730, g19352)
g34076(1) = AND(g33694, g19519)
g33365(1) = AND(g32267, g20994)
g34101(1) = OR(g33693, g33700)
g34231(1) = OR(g33898, g33902)
g34204(1) = OR(g33832, g33833)
g34148(1) = OR(g33758, g19656)
g33353(1) = AND(g32240, g20732)
g34090(1) = OR(g33676, g33680)
g33234(1) = OR(g32039, g32043)
g33374(1) = AND(g32289, g21221)
g34117(1) = AND(g33742, g19755)
g34761(1) = OR(g34679, g34506)
g33933(1) = NAND(g33394, g12491, g12819, g12796)
g34100(1) = OR(g33690, g33697)
g33239(1) = AND(g32117, g19902)
g34166(1) = OR(g33785, g19752)
g34172(1) = OR(g33795, g19914)
g32028(1) = AND(g30569, g29339)
g33227(1) = OR(g32029, g32031)
g34194(1) = OR(g33811, g33815)
g34113(1) = AND(g33734, g19744)
g34743(1) = AND(g8951, g34703)
I31859(1) = OR(g33501, g33502, g33503, g33504)
I31858(1) = OR(g33497, g33498, g33499, g33500)
I31844(1) = OR(g33474, g33475, g33476, g33477)
I31838(1) = OR(g33461, g33462, g33463, g33464)
I31839(1) = OR(g33465, g33466, g33467, g33468)
I31854(1) = OR(g33492, g33493, g33494, g33495)
I31868(1) = OR(g33515, g33516, g33517, g33518)
I31869(1) = OR(g33519, g33520, g33521, g33522)
I31863(1) = OR(g33506, g33507, g33508, g33509)
I31864(1) = OR(g33510, g33511, g33512, g33513)
I31873(1) = OR(g33524, g33525, g33526, g33527)
I31848(1) = OR(g33479, g33480, g33481, g33482)
I31849(1) = OR(g33483, g33484, g33485, g33486)
I31843(1) = OR(g33470, g33471, g33472, g33473)
I31874(1) = OR(g33528, g33529, g33530, g33531)
I31853(1) = OR(g33488, g33489, g33490, g33491)
g30332(1) = NOT(I28597)
g31862(1) = NOT(I29444)
g31863(1) = NOT(I29447)
g33636(1) = NOT(I31463)
g33874(1) = NOT(I31724)
g33935(1) = NOT(I31817)
g34267(1) = OR(g34079, g18728)
g33625(1) = OR(g33373, g18809)
g33624(1) = OR(g33371, g18808)
g34259(1) = OR(g34066, g18679)
g34263(1) = OR(g34078, g18699)
g34023(1) = OR(g33796, g24320)
g33613(1) = OR(g33248, g18649)
g34266(1) = OR(g34076, g18719)
g33623(1) = OR(g33370, g18792)
g33610(1) = OR(g33242, g18616)
g33619(1) = OR(g33359, g18758)
g33614(1) = OR(g33249, g18650)
g33612(1) = OR(g33247, g18633)
g34262(1) = OR(g34075, g18697)
g34268(1) = OR(g34082, g18730)
g34260(1) = OR(g34113, g18680)
g33622(1) = OR(g33366, g18791)
g34849(1) = OR(g34842, g18154)
g33618(1) = OR(g33353, g18757)
g33627(1) = OR(g33376, g18826)
g34269(1) = OR(g34083, g18732)
g34265(1) = OR(g34117, g18711)
g33626(1) = OR(g33374, g18825)
g34264(1) = OR(g34081, g18701)
g34257(1) = OR(g34226, g18674)
g34791(1) = OR(g34771, g18184)
g33620(1) = OR(g33360, g18774)
g34024(1) = OR(g33807, g24331)
g33621(1) = OR(g33365, g18775)
g34261(1) = OR(g34074, g18688)
g33611(1) = OR(g33243, g18632)
g33609(1) = OR(g33239, g18615)
g34258(1) = OR(g34211, g18675)
g33920(1) = NOT(I31786)
g33936(1) = NOT(I31820)
g33682(1) = NOT(I31515)
g33648(4) = NOT(I31482)
g33755(2) = NOT(I31610)
g33845(1) = NOT(I31694)
g33926(1) = NOT(I31796)
g32384(1) = NOT(g31666)
g32382(1) = NOT(g31657)
g33766(5) = NOT(I31619)
I32639(1) = NOT(g34345)
g34132(1) = NOT(g33831)
g33937(4) = NOT(I31823)
g34068(1) = NOT(g33728)
g33120(1) = NOT(I30686)
g33698(1) = NOT(I31539)
g33661(4) = NOT(I31497)
g33888(1) = NOT(g33346)
g32363(1) = NOT(I29891)
g32015(1) = NOT(I29571)
g33931(1) = NOT(I31807)
I29438(1) = NOT(g30610)
I32150(1) = NOT(g33923)
g33658(1) = NOT(g33080)
g33631(4) = NOT(I31459)
g34042(1) = NOT(g33674)
g33875(1) = NOT(I31727)
g34124(1) = NOT(g33819)
g33653(4) = NOT(I31486)
g33917(1) = NOT(I31779)
g33688(1) = NOT(I31523)
g34053(1) = NOT(g33683)
g33456(1) = NOT(I30986)
g33916(1) = NOT(I31776)
g33670(4) = NOT(I31504)
g33335(2) = NOT(I30861)
g33839(1) = NOT(I31686)
g32453(1) = NOT(I29981)
g33800(1) = NOT(I31642)
g33635(1) = NOT(g33436)
g33772(5) = NOT(I31622)
g33641(4) = NOT(I31474)
g33442(1) = NOT(g31937)
g33806(1) = NOT(I31650)
g34049(1) = NOT(g33678)
I29585(1) = NOT(g31655)
g33726(1) = NOT(I31581)
g33791(2) = OR(g33379, g32430)
g32404(2) = NOT(I29936)
I32364(1) = NOT(g34208)
g33750(4) = NOT(I31607)
g33702(1) = NOT(I31545)
g33912(1) = NOT(I31770)
g33691(1) = NOT(I31528)
g33929(1) = NOT(I31803)
g33928(1) = NOT(I31800)
g33827(1) = NOT(I31672)
g34044(1) = NOT(g33675)
g33778(5) = NOT(I31625)
g33932(1) = NOT(I31810)
g34181(1) = NOT(g33913)
g33850(1) = NOT(I31701)
g33716(1) = NOT(I31569)
g34060(1) = NOT(g33704)
g34197(1) = NOT(g33812)
g34070(1) = NOT(g33725)
g30917(1) = NOT(I28897)
g33736(5) = NOT(I31597)
I31535(1) = NOT(g33377)
g33283(2) = OR(g31995, g30318)
g34156(1) = NOT(g33907)
g33708(1) = NOT(I31555)
g33459(1) = NOT(I30995)
g33458(1) = NOT(I30992)
g33918(1) = NOT(I31782)
g33424(1) = NOT(g32415)
g33713(1) = NOT(I31564)
g33705(1) = NOT(I31550)
g33455(1) = NOT(I30983)
g32441(1) = NOT(I29969)
g33665(4) = NOT(I31500)
g33454(1) = NOT(I30980)
g33712(1) = NOT(I31561)
g33637(1) = NOT(I31466)
g33729(1) = NOT(I31586)
g34192(1) = NOT(g33921)
g34062(1) = NOT(g33711)
g33813(1) = NOT(I31659)
g33934(1) = NOT(I31814)
g33761(4) = NOT(I31616)
g33744(5) = NOT(I31604)
g34380(1) = AND(g34158, g20571)
g34811(1) = AND(g14165, g34766)
g33829(1) = AND(g33240, g20164)
g34342(1) = AND(g34103, g19998)
g34393(1) = AND(g34189, g21304)
g34365(1) = AND(g34149, g20451)
g34337(1) = AND(g34095, g19881)
g34171(1) = AND(g33925, g24360)
g34295(1) = AND(g34057, g19370)
g33818(1) = AND(g33236, g20113)
g33735(1) = AND(g33118, g19553)
g34401(1) = AND(g34199, g21383)
g34382(1) = AND(g34167, g20618)
g34284(1) = AND(g34046, g19351)
g34415(1) = AND(g34207, g21458)
g34414(1) = AND(g34206, g21457)
g33727(1) = AND(g33115, g19499)
g33821(1) = AND(g33238, g20153)
g34291(1) = AND(g34055, g19366)
g34173(1) = AND(g33679, g24368)
g34395(1) = AND(g34193, g21336)
g34389(1) = AND(g34170, g20715)
g33731(1) = AND(g33116, g19520)
g34394(1) = AND(g34190, g21305)
g33743(1) = AND(g33119, g19574)
g33803(1) = AND(g33231, g20071)
g34281(1) = AND(g34043, g19276)
g34301(1) = AND(g34064, g19415)
g34120(1) = AND(g33930, g25158)
g34385(1) = AND(g34168, g20642)
g34338(1) = AND(g34099, g19905)
g34867(1) = AND(g34826, g20145)
g34819(1) = OR(g34741, g34684)
g34496(1) = NOR(g34370, g27648)
g34341(1) = AND(g34101, g19952)
g34279(1) = AND(g34231, g19208)
g34410(1) = AND(g34204, g21427)
g34363(1) = AND(g34148, g20389)
g34179(1) = AND(g33686, g24372)
g34334(1) = AND(g34090, g19865)
g33816(1) = AND(g33234, g20096)
g34841(1) = AND(g34761, g20080)
g34116(1) = AND(g33933, g25140)
g34340(1) = AND(g34100, g19950)
g34381(1) = AND(g34166, g20594)
g34390(1) = AND(g34172, g21069)
g34183(1) = AND(g33695, g24385)
g33798(1) = AND(g33227, g20058)
g34396(1) = AND(g34194, g21337)
g33951(1) = OR(g33469, I31838, I31839)
g33957(1) = OR(g33523, I31868, I31869)
g33956(1) = OR(g33514, I31863, I31864)
g33953(1) = OR(g33487, I31848, I31849)
g33952(1) = OR(g33478, I31843, I31844)
g33958(1) = OR(g33532, I31873, I31874)
g33955(1) = OR(g33505, I31858, I31859)
g33954(1) = OR(g33496, I31853, I31854)
g31860(1) = NOT(I29438)
g33945(1) = OR(g32430, g33455)
g33946(1) = OR(g32434, g33456)
g33948(1) = OR(g32442, g33458)
g33949(1) = OR(g32446, g33459)
g34233(1) = OR(g32455, g33951)
g34234(1) = OR(g32520, g33952)
g34235(1) = OR(g32585, g33953)
g34236(1) = OR(g32650, g33954)
g34237(1) = OR(g32715, g33955)
g34238(1) = OR(g32780, g33956)
g34239(1) = OR(g32845, g33957)
g34240(1) = OR(g32910, g33958)
g34441(1) = OR(g34381, g18540)
g34460(1) = OR(g34301, g18677)
g34031(1) = OR(g33735, g18705)
g34452(1) = OR(g34401, g18665)
g34455(1) = OR(g34284, g18668)
g34041(1) = OR(g33829, g18739)
g34448(1) = OR(g34365, g18553)
g34462(1) = OR(g34334, g18685)
g34447(1) = OR(g34363, g18552)
g34446(1) = OR(g34390, g18550)
g34442(1) = OR(g34380, g18542)
g34880(1) = OR(g34867, g18153)
g34451(1) = OR(g34393, g18664)
g34030(1) = OR(g33727, g18704)
g34253(1) = OR(g34171, g24300)
g34033(1) = OR(g33821, g18708)
g34463(1) = OR(g34338, g18686)
g34255(1) = OR(g34120, g24302)
g34464(1) = OR(g34340, g18687)
g34454(1) = OR(g34414, g18667)
g34850(1) = OR(g34841, g18185)
g34458(1) = OR(g34396, g18671)
g34453(1) = OR(g34410, g18666)
g34456(1) = OR(g34395, g18669)
g34038(1) = OR(g33731, g18735)
g34032(1) = OR(g33816, g18706)
g34459(1) = OR(g34415, g18673)
g34040(1) = OR(g33818, g18737)
g34029(1) = OR(g33798, g18703)
g34039(1) = OR(g33743, g18736)
g34444(1) = OR(g34389, g18546)
g34254(1) = OR(g34116, g24301)
g34467(1) = OR(g34341, g18717)
g34256(1) = OR(g34173, g24303)
g34465(1) = OR(g34295, g18712)
g34450(1) = OR(g34281, g18663)
g34468(1) = OR(g34342, g18718)
g34445(1) = OR(g34382, g18548)
g34037(1) = OR(g33803, g18734)
g34443(1) = OR(g34385, g18545)
g34466(1) = OR(g34337, g18716)
g34461(1) = OR(g34291, g18681)
g34449(1) = OR(g34279, g18662)
g34457(1) = OR(g34394, g18670)
g34398(1) = AND(g7684, g34070)
g34188(1) = NOT(g33875)
g34089(1) = AND(g22957, g9104, g33744)
g34229(1) = NOT(g33936)
g34319(1) = AND(g9535, g34156)
g34115(1) = AND(g20516, g9104, g33750)
g34105(1) = AND(g33778, g9104, g18957)
g34080(1) = AND(g22957, g9104, g33750)
g34378(1) = AND(g13095, g34053)
I29441(1) = NOT(g30917)
g33388(1) = NOT(g32382)
g34093(1) = AND(g20114, g33755, g9104)
I32096(1) = NOT(g33641)
I32116(1) = NOT(g33937)
I32093(1) = NOT(g33670)
g34112(1) = AND(g22957, g9104, g33778)
g34358(1) = NOT(I32364)
g34195(1) = NOT(I32150)
g34088(1) = AND(g33736, g9104, g18957)
I31491(1) = NOT(g33283)
I32109(1) = NOT(g33631)
I32119(1) = NOT(g33648)
g34335(1) = AND(g8461, g34197)
I32158(1) = NOT(g33791)
I30989(1) = NOT(g32441)
I32062(1) = NOT(g33653)
I32051(1) = NOT(g33631)
g34086(1) = AND(g20114, g33766, g9104)
I31494(1) = NOT(g33283)
I30971(1) = NOT(g32015)
g34375(1) = AND(g13077, g34049)
g34098(1) = AND(g33744, g9104, g18957)
g34052(1) = NOT(g33635)
g34096(1) = AND(g22957, g9104, g33772)
g33391(1) = NOT(g32384)
I30766(1) = NOT(g32363)
I32056(1) = NOT(g33641)
g32027(1) = NOT(I29585)
I32161(1) = NOT(g33791)
g34092(1) = AND(g33750, g9104, g18957)
I32079(1) = NOT(g33937)
I32106(1) = NOT(g33653)
g34333(1) = AND(g9984, g34192)
g34059(1) = NOT(g33658)
g33696(1) = NOT(I31535)
g34386(1) = AND(g10800, g34060)
I32074(1) = NOT(g33670)
g34298(1) = AND(g8679, g34132)
I32067(1) = NOT(g33661)
g34077(1) = AND(g22957, g9104, g33736)
I31829(1) = NOT(g33454)
g34085(1) = AND(g33761, g9104, g18957)
g34094(1) = NOT(g33772)
I32103(1) = NOT(g33661)
I31361(1) = NOT(g33120)
g34087(1) = AND(g33766, g9104, g18957)
g34329(1) = AND(g14511, g34181)
g34569(1) = NOT(I32639)
I30998(1) = NOT(g32453)
g34371(1) = AND(g7450, g34044)
g34047(1) = NOT(g33637)
I32089(1) = NOT(g33665)
I32071(1) = NOT(g33665)
g34287(1) = AND(g11370, g34124)
g34119(1) = AND(g20516, g9104, g33755)
I32059(1) = NOT(g33648)
g34108(1) = AND(g22957, g9104, g33766)
g34367(1) = AND(g7404, g34042)
g34397(1) = AND(g7673, g34068)
g34091(1) = AND(g22957, g9104, g33761)
g34388(1) = AND(g10802, g34062)
g34097(1) = AND(g33772, g9104, g18957)
g34405(1) = OR(g34183, g25103)
g34182(1) = AND(g33691, g24384)
g34212(1) = AND(g33761, g22689)
g34104(1) = AND(g33916, g23639)
g34133(1) = AND(g33845, g23958)
g34228(1) = AND(g33750, g22942)
g34050(1) = AND(g33772, g22942)
g33899(1) = AND(g32132, g33335)
g34198(1) = AND(g33688, g24491)
g33071(1) = AND(g31591, g32404)
g34225(1) = AND(g33744, g22942)
g34224(1) = AND(g33736, g22670)
g34065(1) = AND(g33813, g23148)
g34219(1) = AND(g33736, g22942)
g34218(1) = AND(g33744, g22670)
g34185(1) = AND(g33702, g24389)
g34215(1) = AND(g33778, g22670)
g34139(1) = AND(g33827, g23314)
g34138(1) = AND(g33929, g23828)
g33110(1) = AND(g32404, g32415)
g34184(1) = AND(g33698, g24388)
g34214(1) = AND(g33772, g22689)
g34114(1) = AND(g33920, g23742)
g34141(1) = AND(g33932, g23828)
g34135(1) = AND(g33926, g23802)
g34106(1) = AND(g33917, g23675)
g34191(1) = AND(g33713, g24404)
g34045(1) = AND(g33766, g22942)
g34140(1) = AND(g33931, g23802)
g34061(1) = AND(g33800, g23076)
g34203(1) = AND(g33726, g24537)
g34196(1) = AND(g33682, g24485)
g34866(1) = AND(g34819, g20106)
g34706(1) = AND(g34496, g10570)
g34102(1) = AND(g33912, g23599)
g33924(1) = AND(g33335, g33346)
g34054(1) = AND(g33778, g22942)
g34180(1) = AND(g33716, g24373)
g34187(1) = AND(g33708, g24397)
g34143(1) = AND(g33934, g23828)
g34217(1) = AND(g33736, g22876)
g34402(1) = OR(g34179, g25084)
g34223(1) = AND(g33744, g22876)
g34178(1) = AND(g33712, g24361)
g34186(1) = AND(g33705, g24396)
g34216(1) = AND(g33778, g22689)
g34856(1) = OR(g34811, g34743)
g34230(1) = AND(g33761, g22942)
g34063(1) = AND(g33806, g23121)
g34137(1) = AND(g33928, g23802)
g34136(1) = AND(g33850, g23293)
g34109(1) = AND(g33918, g23708)
g34213(1) = AND(g33766, g22689)
g34205(1) = AND(g33729, g24541)
g34072(1) = AND(g33839, g24872)
I32185(2) = NAND(g33665, g33661)
I31972(2) = NAND(g33641, g33631)
I31983(2) = NAND(g33653, g33648)
I32202(2) = NAND(g33937, g33670)
g31861(1) = NOT(I29441)
g33533(1) = NOT(I31361)
g33659(1) = NOT(I31491)
g34201(1) = NOT(I32158)
g34881(1) = OR(g34866, g18187)
g34123(1) = NOT(I32062)
I32550(1) = NOT(g34398)
g34134(1) = NOT(I32079)
g34387(1) = NOT(g34188)
g34343(1) = NOT(g34089)
I32601(1) = NOT(g34319)
I32617(1) = NOT(g34333)
g34317(1) = NOT(g34115)
g34323(1) = NOT(g34105)
g34299(1) = NOT(g34080)
I32654(1) = NOT(g34378)
g34316(1) = NOT(g34093)
g34160(1) = NOT(I32119)
g34153(2) = OR(g33899, g33451)
g34145(1) = NOT(I32096)
g34130(1) = NOT(I32071)
g34118(1) = NOT(I32051)
I31477(1) = NOT(g33391)
g34159(1) = NOT(I32116)
g34144(1) = NOT(I32093)
g34336(1) = NOT(g34112)
I30537(1) = NOT(g32027)
I32607(1) = NOT(g34358)
I32274(1) = NOT(g34195)
I31469(1) = NOT(g33388)
g34308(1) = NOT(g34088)
g34202(1) = NOT(I32161)
I32613(1) = NOT(g34329)
g33628(2) = OR(g33071, g32450)
I32621(1) = NOT(g34335)
g33228(2) = NOT(I30766)
g33457(1) = NOT(I30989)
g34151(1) = NOT(I32106)
g34150(1) = NOT(I32103)
g34313(1) = NOT(g34086)
I32284(1) = NOT(g34052)
g33660(1) = NOT(I31494)
g33443(2) = NOT(I30971)
I32651(1) = NOT(g34375)
g34312(1) = NOT(g34098)
g34122(1) = NOT(I32059)
g34142(1) = NOT(I32089)
g34328(1) = NOT(g34096)
g34121(1) = NOT(I32056)
g34325(1) = NOT(g34092)
I32645(1) = NOT(g34367)
g34272(1) = NOT(g34229)
g34737(1) = NOR(g34706, g30003)
g34152(1) = NOT(I32109)
I32547(1) = NOT(g34397)
I31878(1) = NOT(g33696)
I32665(1) = NOT(g34386)
I32594(1) = NOT(g34298)
g34126(1) = NOT(I32067)
g34339(1) = NOT(g34077)
I32297(1) = NOT(g34059)
g33944(1) = NOT(I31829)
g34315(1) = NOT(g34085)
I32699(1) = NOT(g34569)
g34307(1) = NOT(g34087)
g34131(1) = NOT(I32074)
I32671(1) = NOT(g34388)
g33460(1) = NOT(I30998)
I32648(1) = NOT(g34371)
g34275(1) = NOT(g34047)
I32591(1) = NOT(g34287)
g34320(1) = NOT(g34119)
g34327(1) = NOT(g34108)
g34326(1) = NOT(g34091)
g34311(1) = NOT(g34097)
g34482(1) = AND(g34405, g18917)
g34318(1) = OR(g25850, g34063)
g34306(1) = OR(g25782, g34054)
g34305(1) = OR(g25775, g34050)
g34314(1) = OR(g25831, g34061)
g34368(1) = OR(g26274, g34135)
g34274(1) = OR(g27822, g34205)
g34421(1) = OR(g27686, g34198)
g34297(1) = OR(g26858, g34228)
g34417(1) = OR(g27678, g34196)
g34353(1) = OR(g26088, g34114)
g34366(1) = OR(g26257, g34133)
g34399(1) = OR(g34178, g25067)
g34411(1) = OR(g34186, g25142)
g34349(1) = OR(g26019, g34104)
g34377(1) = OR(g26304, g34141)
g34293(1) = OR(g26854, g34224)
g34292(1) = OR(g26853, g34223)
g34376(1) = OR(g26301, g34140)
g34407(1) = OR(g34185, g25124)
g34347(1) = OR(g25986, g34102)
g34288(1) = OR(g26846, g34217)
g34286(1) = OR(g26842, g34216)
g34280(1) = OR(g26833, g34213)
g34331(1) = OR(g27121, g34072)
g34372(1) = OR(g26287, g34137)
g34321(1) = OR(g25866, g34065)
g34369(1) = OR(g26279, g34136)
g34404(1) = OR(g34182, g25102)
g34294(1) = OR(g26855, g34225)
g34303(1) = OR(g25768, g34045)
g34278(1) = OR(g26829, g34212)
g34300(1) = OR(g26864, g34230)
g34416(1) = OR(g34191, g25159)
g34352(1) = OR(g26079, g34109)
g34403(1) = OR(g34180, g25085)
g34478(1) = AND(g34402, g18904)
g34412(1) = OR(g34187, g25143)
g34350(1) = OR(g26048, g34106)
g34909(1) = AND(g34856, g20130)
g34379(1) = OR(g26312, g34143)
g34273(1) = OR(g27765, g34203)
g34290(1) = OR(g26848, g34219)
g34289(1) = OR(g26847, g34218)
g34374(1) = OR(g26294, g34139)
g34406(1) = OR(g34184, g25123)
g34373(1) = OR(g26292, g34138)
g34283(1) = OR(g26839, g34215)
g34282(1) = OR(g26838, g34214)
g34413(1) = AND(g34094, g22670)
I32187(1) = NAND(g33661, I32185)
I32186(1) = NAND(g33665, I32185)
I31984(1) = NAND(g33653, I31983)
I31985(1) = NAND(g33648, I31983)
I31974(1) = NAND(g33631, I31972)
I32204(1) = NAND(g33670, I32202)
I32203(1) = NAND(g33937, I32202)
I31973(1) = NAND(g33641, I31972)
g32975(1) = NOT(I30537)
g33947(1) = OR(g32438, g33457)
g33950(1) = OR(g32450, g33460)
g33959(1) = NOT(I31878)
g34232(1) = OR(g33451, g33944)
g34597(1) = NOT(I32699)
g34911(1) = OR(g34909, g18188)
g34637(1) = OR(g34478, g18694)
g34642(1) = OR(g34482, g18725)
I32243(1) = NOT(g34134)
I32231(1) = NOT(g34123)
g34409(1) = NOT(g34145)
g34470(1) = AND(g7834, g34325)
g34578(1) = AND(g24578, g34308)
g34549(1) = NOT(I32617)
g34408(1) = NOT(g34144)
I32234(1) = NOT(g34126)
g34582(1) = AND(g7764, g34313)
g34420(1) = NOT(g34152)
g34271(1) = NOT(g34160)
I32391(1) = NOT(g34153)
I32237(1) = NOT(g34130)
g34585(1) = AND(g24705, g34316)
I32222(1) = NOT(g34118)
g33645(1) = NOT(I31477)
I31751(1) = NOT(g33228)
g34581(1) = AND(g22864, g34312)
g34392(1) = NOT(g34202)
g34544(1) = NOT(I32613)
g34270(1) = NOT(g34159)
I31748(1) = NOT(g33228)
I32388(1) = NOT(g34153)
I32192(1) = NOT(g33628)
g34277(1) = NOT(I32274)
g34419(1) = NOT(g34151)
g34418(1) = NOT(g34150)
g34058(1) = NOT(g33660)
g34285(1) = NOT(I32284)
g34474(1) = AND(g20083, g34326)
g34502(1) = AND(g26363, g34343)
g34477(1) = AND(g26344, g34328)
g34584(1) = AND(g24653, g34315)
g34400(1) = NOT(g34142)
g34576(1) = NOT(I32654)
I32228(1) = NOT(g34122)
g33638(1) = NOT(I31469)
g34499(1) = AND(g31288, g34339)
I32225(1) = NOT(g34121)
g34491(1) = NOT(I32550)
g34573(1) = NOT(I32645)
I32240(1) = NOT(g34131)
I32195(1) = NOT(g33628)
g34498(1) = AND(g13888, g34336)
g34844(1) = NOT(g34737)
g34540(1) = NOT(I32607)
g34571(1) = AND(g27225, g34299)
g34586(1) = AND(g11025, g34317)
g34490(1) = NOT(I32547)
g34296(1) = NOT(I32297)
g34588(1) = AND(g26082, g34323)
g34531(1) = NOT(I32594)
g34587(1) = NOT(I32671)
g34577(1) = AND(g24577, g34307)
g34580(1) = AND(g29539, g34311)
g34530(1) = NOT(I32591)
g34575(1) = NOT(I32651)
g34553(1) = NOT(I32621)
g34536(1) = NOT(I32601)
g34475(1) = AND(g27450, g34327)
g34574(1) = NOT(I32648)
g34583(1) = NOT(I32665)
g34533(1) = AND(g34318, g19731)
g34529(1) = AND(g34306, g19634)
g34528(1) = AND(g34305, g19617)
g34532(1) = AND(g34314, g19710)
g34561(1) = AND(g34368, g17410)
g34495(1) = AND(g34274, g19365)
g34489(1) = AND(g34421, g19068)
g34525(1) = AND(g34297, g19528)
g34488(1) = AND(g34417, g18988)
g34558(1) = AND(g34353, g20578)
g34494(1) = OR(g26849, g34413)
g34560(1) = AND(g34366, g17366)
g34476(1) = AND(g34399, g18891)
g34485(1) = AND(g34411, g18952)
g34555(1) = AND(g34349, g20512)
g34567(1) = AND(g34377, g17491)
g34519(1) = AND(g34293, g19504)
g34518(1) = AND(g34292, g19503)
g33677(1) = AND(g33443, g31937)
g34566(1) = AND(g34376, g17489)
g34484(1) = AND(g34407, g18939)
g34554(1) = AND(g34347, g20495)
g34515(1) = AND(g34288, g19491)
g34514(1) = AND(g34286, g19480)
g34507(1) = AND(g34280, g19454)
g34541(1) = AND(g34331, g20087)
g34563(1) = AND(g34372, g17465)
g34534(1) = AND(g34321, g19743)
g34562(1) = AND(g34369, g17411)
g34481(1) = AND(g34404, g18916)
g34572(1) = AND(g34387, g33326)
g34520(1) = AND(g34294, g19505)
g34497(1) = AND(g34275, g33072)
g34527(1) = AND(g34303, g19603)
g34503(1) = AND(g34278, g19437)
g34526(1) = AND(g34300, g19569)
g33657(1) = AND(g30991, g33443)
g34487(1) = AND(g34416, g18983)
g34557(1) = AND(g34352, g20555)
g34479(1) = AND(g34403, g18905)
g34486(1) = AND(g34412, g18953)
g34556(1) = AND(g34350, g20537)
g34568(1) = AND(g34379, g17512)
g34493(1) = AND(g34273, g19360)
g34517(1) = AND(g34290, g19493)
g34516(1) = AND(g34289, g19492)
g34565(1) = AND(g34374, g17471)
g34492(1) = AND(g34272, g33430)
g34483(1) = AND(g34406, g18938)
g34564(1) = AND(g34373, g17466)
g34509(1) = AND(g34283, g19473)
g34508(1) = AND(g34282, g19472)
g34056(2) = NAND(I31984, I31985)
g34051(2) = NAND(I31973, I31974)
g34220(2) = NAND(I32186, I32187)
g34227(2) = NAND(I32203, I32204)
g33894(1) = NOT(I31748)
g34221(1) = NOT(I32192)
g34383(1) = NOT(I32388)
g34617(1) = OR(g34526, g18579)
g34646(1) = OR(g34557, g18803)
g34609(1) = OR(g34503, g18563)
g34645(1) = OR(g34556, g18786)
g34644(1) = OR(g34555, g18769)
g34627(1) = OR(g34534, g18644)
g34636(1) = OR(g34476, g18693)
g34643(1) = OR(g34554, g18752)
g34625(1) = OR(g34532, g18610)
g34610(1) = OR(g34507, g18564)
g34638(1) = OR(g34484, g18721)
g34622(1) = OR(g34520, g18584)
g34605(1) = OR(g34566, g15077)
g34598(1) = OR(g34541, g18136)
g34647(1) = OR(g34558, g18820)
g34603(1) = OR(g34561, g15075)
g34611(1) = OR(g34508, g18565)
g34626(1) = OR(g34533, g18627)
g34628(1) = OR(g34493, g18653)
g34634(1) = OR(g34483, g18691)
g34624(1) = OR(g34509, g18592)
g34639(1) = OR(g34486, g18722)
g34641(1) = OR(g34479, g18724)
g34629(1) = OR(g34495, g18654)
g34640(1) = OR(g34487, g18723)
g34615(1) = OR(g34516, g18576)
g34604(1) = OR(g34563, g15076)
g34602(1) = OR(g34489, g18269)
g34631(1) = OR(g34562, g15118)
g34613(1) = OR(g34515, g18567)
g34616(1) = OR(g34519, g18577)
g34632(1) = OR(g34565, g15119)
g34606(1) = OR(g34564, g15080)
g34621(1) = OR(g34517, g18583)
g34633(1) = OR(g34481, g18690)
g34635(1) = OR(g34485, g18692)
g34601(1) = OR(g34488, g18211)
g34607(1) = OR(g34567, g15081)
g34620(1) = OR(g34529, g18582)
g34619(1) = OR(g34528, g18581)
g34614(1) = OR(g34518, g18568)
g34608(1) = OR(g34568, g15082)
g34618(1) = OR(g34527, g18580)
g34630(1) = OR(g34560, g15117)
g34612(1) = OR(g34514, g18566)
g34623(1) = OR(g34525, g18585)
g34248(1) = NOT(I32243)
g34511(1) = NOT(g34419)
I32800(1) = NOT(g34582)
g34505(1) = NOT(g34409)
I32815(1) = NOT(g34470)
I32791(1) = NOT(g34578)
g34504(1) = NOT(g34408)
g34245(1) = NOT(I32234)
g34512(1) = NOT(g34420)
I32806(1) = NOT(g34585)
g34244(1) = NOT(I32231)
g33895(1) = NOT(I31751)
I32820(1) = NOT(g34474)
I32797(1) = NOT(g34581)
I32788(1) = NOT(g34577)
g34384(1) = NOT(I32391)
g34708(1) = OR(g33381, g34572)
g34241(1) = NOT(I32222)
g34276(1) = NOT(g34058)
I32846(1) = NOT(g34502)
g34649(1) = OR(g33111, g34492)
g34570(1) = NOT(g34392)
I32827(1) = NOT(g34477)
I32803(1) = NOT(g34584)
I32809(1) = NOT(g34586)
g34501(1) = NOT(g34400)
g34127(2) = OR(g33657, g32438)
I32782(1) = NOT(g34571)
I32476(1) = NOT(g34277)
I32843(1) = NOT(g34499)
I32824(1) = NOT(g34475)
g34243(1) = NOT(I32228)
g34521(1) = NOT(g34270)
g34247(1) = NOT(I32240)
g34510(1) = NOT(g34418)
I32525(1) = NOT(g34285)
g34246(1) = NOT(I32237)
I32837(1) = NOT(g34498)
g34242(1) = NOT(I32225)
I32170(1) = NOT(g33638)
I32855(1) = NOT(g34540)
g34657(1) = OR(g33114, g34497)
I32535(1) = NOT(g34296)
I32794(1) = NOT(g34580)
I32173(1) = NOT(g33645)
I32812(1) = NOT(g34588)
g34222(1) = NOT(I32195)
g34522(1) = NOT(g34271)
g34710(1) = AND(g34553, g20903)
g34681(1) = AND(g34491, g19438)
g34696(1) = AND(g34531, g20004)
g34709(1) = AND(g34549, g17242)
g34678(1) = AND(g34490, g19431)
g34686(1) = AND(g34494, g19494)
g34665(1) = AND(g34583, g19067)
g34701(1) = AND(g34536, g20179)
g34661(1) = AND(g34575, g18907)
g34658(1) = AND(g34574, g18896)
g34707(1) = AND(g34544, g20579)
g34876(1) = AND(g34844, g20534)
g34655(1) = AND(g34573, g18885)
g34694(1) = AND(g34530, g19885)
g34666(1) = AND(g34587, g19144)
g34662(1) = AND(g34576, g18931)
I32431(2) = NAND(g34056, g34051)
I32439(2) = NAND(g34227, g34220)
g34435(1) = NOT(I32476)
g34733(1) = OR(g34678, g18651)
g34882(1) = OR(g34876, g18659)
g34727(1) = OR(g34655, g18213)
g34729(1) = OR(g34666, g18270)
g34730(1) = OR(g34658, g18271)
g34726(1) = OR(g34665, g18212)
g34719(1) = OR(g34701, g18133)
g34721(1) = OR(g34696, g18135)
g34720(1) = OR(g34694, g18134)
g34731(1) = OR(g34662, g18272)
g34734(1) = OR(g34681, g18652)
g34732(1) = OR(g34686, g18593)
g34722(1) = OR(g34707, g18137)
g34728(1) = OR(g34661, g18214)
g34723(1) = OR(g34710, g18139)
g34735(1) = OR(g34709, g15116)
I32763(1) = NOT(g34511)
g34672(1) = NOT(I32800)
I32470(1) = NOT(g34247)
I32878(1) = NOT(g34501)
I32458(1) = NOT(g34243)
I32455(1) = NOT(g34242)
I32467(1) = NOT(g34246)
I32904(1) = NOT(g34708)
g34423(1) = NOT(g34222)
I32446(1) = NOT(g34127)
I32770(1) = NOT(g34505)
g34680(1) = NOT(I32820)
g34472(1) = NOT(I32525)
I32464(1) = NOT(g34245)
g34669(1) = NOT(I32791)
g34668(1) = NOT(I32788)
g34559(1) = NOT(g34384)
I32871(1) = NOT(g34521)
g34480(1) = NOT(I32535)
I32452(1) = NOT(g34241)
I32929(1) = NOT(g34649)
g34675(1) = NOT(I32809)
I32449(1) = NOT(g34127)
g34664(1) = NOT(I32782)
g34200(1) = NOT(g33895)
g34674(1) = NOT(I32806)
g34692(1) = NOT(I32846)
g34683(1) = NOT(I32827)
I32775(1) = NOT(g34512)
I32935(1) = NOT(g34657)
I32461(1) = NOT(g34244)
I32473(1) = NOT(g34248)
g34682(1) = NOT(I32824)
I32752(1) = NOT(g34510)
g34210(1) = NOT(I32173)
g34699(1) = NOT(I32855)
g34209(1) = NOT(I32170)
I32874(1) = NOT(g34504)
g34671(1) = NOT(I32797)
g34689(1) = NOT(I32837)
g34670(1) = NOT(I32794)
g34677(1) = NOT(I32815)
g34676(1) = NOT(I32812)
I32766(1) = NOT(g34522)
g34673(1) = NOT(I32803)
g34691(1) = NOT(I32843)
g34500(1) = AND(g34276, g30568)
g34715(1) = AND(g34570, g33375)
I32440(1) = NAND(g34227, I32439)
I32441(1) = NAND(g34220, I32439)
I32433(1) = NAND(g34051, I32431)
I32432(1) = NAND(g34056, I32431)
g34425(1) = NOT(I32446)
I32976(1) = NOT(g34699)
g34433(1) = NOT(I32470)
g34716(1) = NOT(I32878)
g34429(1) = NOT(I32458)
g34428(1) = NOT(I32455)
I32840(1) = NOT(g34480)
g34656(1) = NOT(I32770)
g34432(1) = NOT(I32467)
g34736(1) = NOT(I32904)
g34471(1) = NOT(g34423)
g34430(1) = NOT(I32461)
I32834(1) = NOT(g34472)
g34713(1) = NOT(I32871)
I32309(1) = NOT(g34210)
g34653(1) = NOT(I32763)
g34759(1) = NOT(I32935)
g34755(1) = NOT(I32929)
g34781(1) = OR(g33431, g34715)
g34434(1) = NOT(I32473)
g34426(1) = NOT(I32449)
g34648(1) = NOT(I32752)
g34431(1) = NOT(I32464)
g34663(1) = OR(g32028, g34500)
g34427(1) = NOT(I32452)
I32305(1) = NOT(g34209)
g34659(1) = NOT(I32775)
g34714(1) = NOT(I32874)
g34654(1) = NOT(I32766)
g34391(1) = NOT(g34200)
g34711(1) = NOT(g34559)
g34765(1) = AND(g34692, g20057)
g34753(1) = AND(g34676, g19586)
g34764(1) = AND(g34691, g20009)
g34752(1) = AND(g34675, g19544)
g34748(1) = AND(g34672, g19529)
g34745(1) = AND(g34669, g19482)
g34758(1) = AND(g34683, g19657)
g34744(1) = AND(g34668, g19481)
g34754(1) = AND(g34677, g19602)
g34763(1) = AND(g34689, g19915)
g34740(1) = AND(g34664, g19414)
g34747(1) = AND(g34671, g19527)
g34751(1) = AND(g34674, g19543)
g34746(1) = AND(g34670, g19526)
g34750(1) = AND(g34673, g19542)
g34757(1) = AND(g34682, g19635)
g34756(1) = AND(g34680, g19618)
g34424(2) = NAND(I32440, I32441)
g34422(2) = NAND(I32432, I32433)
g34807(1) = OR(g34764, g18596)
g34806(1) = OR(g34763, g18595)
g34800(1) = OR(g34752, g18586)
g34795(1) = OR(g34753, g18572)
g34798(1) = OR(g34754, g18575)
g34792(1) = OR(g34750, g18569)
g34804(1) = OR(g34740, g18591)
g34801(1) = OR(g34756, g18588)
g34808(1) = OR(g34765, g18599)
g34797(1) = OR(g34747, g18574)
g34796(1) = OR(g34745, g18573)
g34794(1) = OR(g34746, g18571)
g34803(1) = OR(g34758, g18590)
g34802(1) = OR(g34757, g18589)
g34799(1) = OR(g34751, g18578)
g34793(1) = OR(g34744, g18570)
g34805(1) = OR(g34748, g18594)
g34778(2) = NOT(I32976)
I32988(1) = NOT(g34755)
g34690(1) = NOT(I32840)
g34302(1) = NOT(I32305)
I32953(1) = NOT(g34656)
I32967(1) = NOT(g34648)
I32684(1) = NOT(g34430)
I33020(1) = NOT(g34781)
I32693(1) = NOT(g34433)
I32675(1) = NOT(g34427)
I32690(1) = NOT(g34432)
g34688(1) = NOT(I32834)
g34304(1) = NOT(I32309)
I32681(1) = NOT(g34429)
I32696(1) = NOT(g34434)
I32960(1) = NOT(g34653)
g34473(1) = NOT(g34426)
I32970(1) = NOT(g34716)
I32938(1) = NOT(g34663)
I32956(1) = NOT(g34654)
I32947(1) = NOT(g34659)
I32687(1) = NOT(g34431)
I32985(1) = NOT(g34736)
I32973(1) = NOT(g34714)
I32678(1) = NOT(g34428)
I32991(1) = NOT(g34759)
I32659(1) = NOT(g34391)
I32950(1) = NOT(g34713)
g34782(1) = AND(g34711, g33888)
g34667(1) = AND(g34471, g33424)
I32516(2) = NAND(g34424, g34422)
g34593(1) = NOT(I32687)
g34787(1) = NOT(I32991)
g34596(1) = NOT(I32696)
g34592(1) = NOT(I32684)
g34589(1) = NOT(I32675)
g34591(1) = NOT(I32681)
g34595(1) = NOT(I32693)
g34785(1) = NOT(I32985)
g34590(1) = NOT(I32678)
g34594(1) = NOT(I32690)
g34786(1) = NOT(I32988)
I32881(1) = NOT(g34688)
g34775(1) = NOT(I32967)
I32884(1) = NOT(g34690)
I32479(1) = NOT(g34302)
g34783(1) = OR(g33110, g34667)
g34810(1) = NOT(I33020)
g34772(1) = NOT(I32960)
I32482(1) = NOT(g34304)
g34769(1) = NOT(I32953)
g34776(1) = NOT(I32970)
g34579(1) = NOT(I32659)
g34767(1) = NOT(I32947)
g34760(1) = NOT(I32938)
g34770(1) = NOT(I32956)
g34777(1) = NOT(I32973)
I33056(1) = NOT(g34778)
g34768(1) = NOT(I32950)
g34660(1) = NOT(g34473)
g34843(1) = OR(g33924, g34782)
I33053(1) = NOT(g34778)
I32517(1) = NAND(g34424, I32516)
I32518(1) = NAND(g34422, I32516)
g34436(1) = NOT(I32479)
g34437(1) = NOT(I32482)
g34839(1) = NOT(I33053)
g34717(1) = NOT(I32881)
g34718(1) = NOT(I32884)
I33044(1) = NOT(g34775)
I33024(1) = NOT(g34783)
I33070(1) = NOT(g34810)
I33037(1) = NOT(g34770)
I33030(1) = NOT(g34768)
I33050(1) = NOT(g34777)
g34840(1) = NOT(I33056)
I33041(1) = NOT(g34772)
I32868(1) = NOT(g34579)
I33034(1) = NOT(g34769)
I33027(1) = NOT(g34767)
I33047(1) = NOT(g34776)
I32997(1) = NOT(g34760)
I33075(1) = NOT(g34843)
g34738(1) = AND(g34660, g33442)
g34469(2) = NAND(I32517, I32518)
g34789(1) = NOT(I32997)
g34848(1) = NOT(I33070)
g34712(1) = NOT(I32868)
g34812(1) = NOT(I33024)
g34823(2) = NOT(I33037)
g34816(2) = NOT(I33030)
g34830(2) = NOT(I33044)
g34836(2) = NOT(I33050)
g34864(1) = NOT(g34840)
g34851(1) = NOT(I33075)
g34813(2) = NOT(I33027)
g34833(2) = NOT(I33047)
g34809(1) = OR(g33677, g34738)
g34820(2) = NOT(I33034)
g34827(2) = NOT(I33041)
I32756(2) = NAND(g34469, g25779)
I32909(1) = NOT(g34712)
I33067(1) = NOT(g34812)
I33109(1) = NOT(g34851)
g34910(1) = NOT(g34864)
I33079(1) = NOT(g34809)
g34857(1) = AND(g16540, g34813)
g34869(1) = AND(g34816, g19869)
g34868(1) = AND(g34813, g19866)
g34865(1) = AND(g16540, g34836)
g34875(1) = AND(g34836, g20073)
g34874(1) = AND(g34833, g20060)
g34861(1) = AND(g16540, g34827)
g34871(1) = AND(g34823, g19908)
g34859(1) = AND(g16540, g34820)
g34858(1) = AND(g16540, g34816)
g34860(1) = AND(g16540, g34823)
g34870(1) = AND(g34820, g19882)
g34863(1) = AND(g16540, g34833)
g34873(1) = AND(g34830, g20046)
g34862(1) = AND(g16540, g34830)
g34872(1) = AND(g34827, g19954)
I32757(1) = NAND(g34469, I32756)
I32758(1) = NAND(g25779, I32756)
g34847(1) = NOT(I33067)
g34879(1) = NOT(I33109)
g34903(2) = OR(g34859, g21690)
g34906(2) = OR(g34857, g21694)
g34884(2) = OR(g34858, g21666)
g34894(2) = OR(g34862, g21678)
g34900(2) = OR(g34860, g21686)
g34739(1) = NOT(I32909)
I33182(1) = NOT(g34910)
g34897(2) = OR(g34861, g21682)
g34855(1) = NOT(I33079)
g34650(2) = NAND(I32757, I32758)
g34890(2) = OR(g34863, g21674)
g34887(2) = OR(g34865, g21670)
I33146(1) = NOT(g34903)
I33167(1) = NOT(g34890)
g34930(1) = NOT(I33182)
I33164(1) = NOT(g34894)
I33106(1) = NOT(g34855)
I33149(1) = NOT(g34900)
I33131(1) = NOT(g34906)
I33143(1) = NOT(g34903)
I33137(1) = NOT(g34884)
I32921(1) = NOT(g34650)
I33134(1) = NOT(g34906)
I33155(1) = NOT(g34897)
I33152(1) = NOT(g34900)
I32994(1) = NOT(g34739)
I33173(1) = NOT(g34887)
I33170(1) = NOT(g34890)
I33161(1) = NOT(g34894)
I33158(1) = NOT(g34897)
I32963(1) = NOT(g34650)
I33140(1) = NOT(g34884)
I33176(1) = NOT(g34887)
g34788(1) = NOT(I32994)
g34913(1) = NOT(I33131)
g34915(1) = NOT(I33137)
g34917(1) = NOT(I33143)
g34919(1) = NOT(I33149)
g34921(1) = NOT(I33155)
g34923(1) = NOT(I33161)
g34925(1) = NOT(I33167)
g34927(1) = NOT(I33173)
g34878(1) = NOT(I33106)
g34914(1) = NOT(I33134)
I33197(1) = NOT(g34930)
g34924(1) = NOT(I33164)
g34918(1) = NOT(I33146)
g34749(1) = NOT(I32921)
g34922(1) = NOT(I33158)
g34920(1) = NOT(I33152)
g34926(1) = NOT(I33170)
g34773(1) = NOT(I32963)
g34916(1) = NOT(I33140)
g34928(1) = NOT(I33176)
g34933(1) = NOT(g34916)
g34932(1) = NOT(g34914)
g34943(1) = NOT(I33197)
I32982(1) = NOT(g34749)
g34939(1) = NOT(g34922)
g34938(1) = NOT(g34920)
g34941(1) = NOT(g34926)
g34845(1) = NOT(g34773)
g34934(1) = NOT(g34918)
g34940(1) = NOT(g34924)
g34942(1) = NOT(g34928)
g34945(1) = NOT(g34933)
g34944(1) = NOT(g34932)
I33210(1) = NOT(g34943)
g34852(2) = NOT(g34845)
g34947(1) = NOT(g34938)
g34951(1) = NOT(g34941)
g34946(1) = NOT(g34934)
g34950(1) = NOT(g34940)
g34784(1) = NOT(I32982)
g34952(1) = NOT(g34942)
g34949(1) = NOT(g34939)
g34954(1) = NOT(I33210)
I33119(1) = NOT(g34852)
g34883(1) = NOT(g34852)
I33064(1) = NOT(g34784)
g34961(1) = AND(g34944, g23019)
g34967(1) = AND(g34951, g23189)
g34966(1) = AND(g34950, g23170)
g34963(1) = AND(g34946, g23041)
g34962(1) = AND(g34945, g23020)
g34968(1) = AND(g34952, g23203)
g34965(1) = AND(g34949, g23084)
g34964(1) = AND(g34947, g23060)
g34970(1) = OR(g34868, g34961)
g34846(1) = NOT(I33064)
g34893(1) = NOT(I33119)
g34978(1) = OR(g34874, g34967)
g34974(1) = OR(g34870, g34963)
g34971(1) = OR(g34869, g34962)
g34977(1) = OR(g34873, g34966)
g34976(1) = OR(g34872, g34965)
I33214(1) = NOT(g34954)
g34975(1) = OR(g34871, g34964)
g34979(1) = OR(g34875, g34968)
g34912(1) = NOR(g34883, g20277, g20242, g21370)
g34956(1) = NOT(I33214)
I33246(1) = NOT(g34970)
I33103(1) = NOT(g34846)
I33267(1) = NOT(g34979)
I33264(1) = NOT(g34978)
I33255(1) = NOT(g34975)
I33179(1) = NOT(g34893)
I33252(1) = NOT(g34974)
I33249(1) = NOT(g34971)
I33261(1) = NOT(g34977)
I33258(1) = NOT(g34976)
g34931(1) = OR(g2984, g34912)
g34877(1) = NOT(I33103)
g34989(1) = NOT(I33267)
g34988(1) = NOT(I33264)
g34986(1) = NOT(I33258)
g34985(1) = NOT(I33255)
g34984(1) = NOT(I33252)
g34987(1) = NOT(I33261)
g34929(1) = NOT(I33179)
g34982(1) = NOT(I33246)
g34955(1) = AND(g34931, g34320)
g34983(1) = NOT(I33249)
I33285(1) = NOT(g34988)
I33218(1) = NOT(g34955)
I33282(1) = NOT(g34987)
I33279(1) = NOT(g34986)
I33189(1) = NOT(g34929)
I33273(1) = NOT(g34984)
I33270(1) = NOT(g34982)
I33291(1) = NOT(g34983)
I33288(1) = NOT(g34989)
I33276(1) = NOT(g34985)
g34993(1) = NOT(I33279)
g34997(1) = NOT(I33291)
g34996(1) = NOT(I33288)
g34991(1) = NOT(I33273)
g34990(1) = NOT(I33270)
g34992(1) = NOT(I33276)
g34995(1) = NOT(I33285)
g34994(1) = NOT(I33282)
g34960(1) = NOT(I33218)
g34935(2) = NOT(I33189)
g34969(1) = AND(g34960, g19570)
g34953(1) = AND(g34935, g19957)
g34948(1) = AND(g16540, g34935)
g34980(1) = OR(g34969, g18587)
g34957(2) = OR(g34948, g21662)
I33235(1) = NOT(g34957)
I33232(1) = NOT(g34957)
g34972(1) = NOT(I33232)
g34973(1) = NOT(I33235)
g34981(1) = NOT(g34973)
g34998(1) = NOT(g34981)
g34999(1) = AND(g34998, g23085)
g35000(1) = OR(g34953, g34999)
I33297(1) = NOT(g35000)
g35001(1) = NOT(I33297)
I33300(1) = NOT(g35001)
g35002(1) = NOT(I33300)
