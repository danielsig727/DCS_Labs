# INPUT 54
# OUTPUT 42
# NOT 254
# AND 94
# OR 17
# NAND 28
INPUT(G1)
INPUT(G2)
INPUT(G3)
INPUT(G4)
INPUT(G5)
INPUT(G6)
INPUT(G8)
INPUT(G9)
INPUT(G10)
INPUT(G11)
INPUT(G12)
INPUT(G13)
INPUT(G14)
INPUT(G15)
INPUT(G16)
INPUT(G17)
INPUT(G18)
INPUT(G19)
INPUT(G20)
INPUT(G21)
INPUT(G22)
INPUT(G23)
INPUT(G24)
INPUT(G25)
INPUT(G26)
INPUT(G27)
INPUT(G28)
INPUT(G29)
INPUT(G30)
INPUT(G31)
INPUT(G32)
INPUT(G33)
INPUT(G34)
INPUT(G35)
INPUT(G36)
INPUT(G64)
INPUT(G65)
INPUT(G66)
INPUT(G67)
INPUT(G68)
INPUT(G69)
INPUT(G70)
INPUT(G71)
INPUT(G72)
INPUT(G73)
INPUT(G74)
INPUT(G75)
INPUT(G76)
INPUT(G77)
INPUT(G78)
INPUT(G79)
INPUT(G80)
INPUT(G81)
INPUT(G82)
OUTPUT(G103BF)
OUTPUT(G104BF)
OUTPUT(G105BF)
OUTPUT(G106BF)
OUTPUT(G107)
OUTPUT(G83)
OUTPUT(G84)
OUTPUT(G85)
OUTPUT(G86BF)
OUTPUT(G87BF)
OUTPUT(G88BF)
OUTPUT(G89BF)
OUTPUT(G90)
OUTPUT(G91)
OUTPUT(G92)
OUTPUT(G94)
OUTPUT(G95BF)
OUTPUT(G96BF)
OUTPUT(G97BF)
OUTPUT(G98BF)
OUTPUT(G99BF)
OUTPUT(G100BF)
OUTPUT(G101BF)
OUTPUT(G380)
OUTPUT(G262)
OUTPUT(G394)
OUTPUT(G250)
OUTPUT(G122)
OUTPUT(G133)
OUTPUT(G138)
OUTPUT(G139)
OUTPUT(G140)
OUTPUT(G141)
OUTPUT(G142)
OUTPUT(G125)
OUTPUT(G126)
OUTPUT(G127)
OUTPUT(G128)
OUTPUT(G129)
OUTPUT(G130)
OUTPUT(G131)
OUTPUT(G132)
I633(1) = NOT(G1)
G366(1) = NOT(G2)
G379(1) = NOT(G3)
I643(1) = NOT(G4)
I646(1) = NOT(G5)
I649(1) = NOT(G6)
I652(1) = NOT(G8)
I655(1) = NOT(G9)
I660(1) = NOT(G10)
I680(1) = NOT(G11)
I684(1) = NOT(G12)
I687(1) = NOT(G13)
I165(1) = NOT(G27)
II178(1) = NOT(G29)
I169(1) = NOT(G70)
I172(1) = NOT(G71)
I175(1) = NOT(G72)
I178(1) = NOT(G80)
I181(1) = NOT(G73)
I184(1) = NOT(G81)
I187(1) = NOT(G74)
I190(1) = NOT(G82)
I193(1) = NOT(G75)
I196(1) = NOT(G68)
I199(1) = NOT(G76)
I202(1) = NOT(G69)
I205(1) = NOT(G77)
I208(1) = NOT(G78)
I211(1) = NOT(G79)
G91(1) = NOT(I165)
G94(1) = NOT(II178)
G113(1) = NOT(I169)
G115(1) = NOT(I172)
G117(1) = NOT(I175)
G219(1) = NOT(I178)
G119(1) = NOT(I181)
G221(1) = NOT(I184)
G121(1) = NOT(I187)
G223(1) = NOT(I190)
G209(1) = NOT(I193)
G109(1) = NOT(I196)
G211(1) = NOT(I199)
G111(1) = NOT(I202)
G213(1) = NOT(I205)
G215(1) = NOT(I208)
G217(1) = NOT(I211)
G352(1) = NOT(I633)
G360(1) = NOT(I643)
G361(1) = NOT(I646)
G362(1) = NOT(I649)
G363(1) = NOT(I652)
G364(1) = NOT(I655)
G367(1) = NOT(I660)
G386(1) = NOT(I680)
G388(1) = NOT(I684)
G389(1) = NOT(I687)
G110(1) = NOT(G360)
G114(1) = NOT(G360)
G118(1) = NOT(G360)
G216(1) = NOT(G360)
G218(1) = NOT(G360)
G220(1) = NOT(G360)
G222(1) = NOT(G360)
G365(1) = NOT(G364)
G368(1) = NOT(G367)
G387(1) = NOT(G386)
G225(1) = NOT(G388)
G390(1) = NOT(G389)
G289(1) = AND(G386, G388, G389)
I356(1) = NOT(G289)
G324(1) = AND(G110, G111)
G338(1) = AND(G114, G115)
G344(1) = AND(G118, G119)
G312(1) = AND(G216, G217)
G315(1) = AND(G218, G219)
G318(1) = AND(G220, G221)
G321(1) = AND(G222, G223)
G231(1) = AND(G379, G387)
G232(1) = AND(G379, G387)
G233(1) = AND(G379, G387)
G234(1) = AND(G379, G387)
G247(1) = AND(G379, G365, G368, G390)
G248(1) = AND(G379, G365, G367, G390)
G263(1) = AND(G379, G364, G368, G390)
G264(1) = AND(G379, G364, G367, G390)
I254(1) = NOT(G324)
I257(1) = NOT(G324)
I260(1) = NOT(G338)
I263(1) = NOT(G338)
I266(1) = NOT(G344)
I269(1) = NOT(G344)
I272(1) = NOT(G312)
I275(1) = NOT(G315)
I278(1) = NOT(G318)
I281(1) = NOT(G321)
G143(1) = NOT(I356)
G281(1) = OR(G232, G248, G65)
G283(1) = OR(G234, G67, G264)
G166(1) = NOT(I254)
G325(1) = NOT(I257)
G194(1) = NOT(I260)
G339(1) = NOT(I263)
G202(1) = NOT(I266)
G345(1) = NOT(I269)
G313(1) = NOT(I272)
G316(1) = NOT(I275)
G319(1) = NOT(I278)
G322(1) = NOT(I281)
I303(1) = NOT(G143)
I299(1) = NOT(G281)
I313(1) = NOT(G283)
G107(1) = AND(G313, G18)
G83(1) = AND(G316, G19)
G84(1) = AND(G319, G20)
G85(1) = AND(G322, G21)
I287(1) = NOT(G166)
I291(1) = NOT(G194)
I295(1) = NOT(G202)
G350(1) = NOT(I303)
G100(1) = AND(G325, G35)
G98(1) = AND(G339, G33)
G96(1) = AND(G345, G31)
I301(1) = NOT(I299)
I315(1) = NOT(I313)
I300(1) = NAND(G281, I299)
I314(1) = NAND(G283, I313)
G92(1) = AND(G350, G28)
G96BF(1) = NOT(G96)
G98BF(1) = NOT(G98)
G100BF(1) = NOT(G100)
G381(1) = NOT(I287)
G375(1) = NOT(I291)
G371(1) = NOT(I295)
G135(1) = NAND(I300, I301)
G137(1) = NAND(I314, I315)
G382(1) = NOT(G381)
G376(1) = NOT(G375)
G372(1) = NOT(G371)
I321(1) = NOT(G135)
I324(1) = NOT(G137)
G329(1) = NOT(I321)
G333(1) = NOT(I324)
G87(1) = AND(G329, G23)
G89(1) = AND(G333, G25)
G87BF(1) = NOT(G87)
G89BF(1) = NOT(G89)
I406(1) = NOT(G87)
I422(1) = NOT(G89)
G173(1) = NOT(I406)
G183(1) = NOT(I422)
I335(1) = NOT(G173)
I338(1) = NOT(G183)
G174(1) = NOT(I335)
G184(1) = NOT(I338)
I341(1) = NOT(G174)
G359(1) = NOT(G184)
G355(1) = NOT(I341)
G108(1) = NOT(G359)
G214(1) = NAND(G379, G359)
G356(1) = NOT(G355)
G293(1) = AND(G108, G109)
G309(1) = AND(G214, G215)
G116(1) = NOT(G356)
I354(1) = NOT(G293)
I357(1) = NOT(G293)
I360(1) = NOT(G309)
I363(1) = NOT(G309)
G210(1) = NAND(G379, G356)
G146(1) = NOT(I354)
G294(1) = NOT(I357)
G162(1) = NOT(I360)
G310(1) = NOT(I363)
G341(1) = AND(G116, G117)
G303(1) = AND(G210, G211)
I366(1) = NOT(G341)
I369(1) = NOT(G341)
I372(1) = NOT(G303)
I375(1) = NOT(G303)
I378(1) = NOT(G146)
I382(1) = NOT(G162)
G101(1) = AND(G294, G36)
G106(1) = AND(G310, G17)
G106BF(1) = NOT(G106)
G101BF(1) = NOT(G101)
G198(1) = NOT(I366)
G342(1) = NOT(I369)
G154(1) = NOT(I372)
G304(1) = NOT(I375)
G383(1) = NOT(I378)
G396(1) = NOT(I382)
G250(1) = AND(G366, G396)
I386(1) = NOT(G198)
I390(1) = NOT(G154)
G384(1) = NOT(G383)
G397(1) = NOT(G396)
G97(1) = AND(G342, G32)
G104(1) = AND(G304, G15)
G278(1) = AND(G366, G396)
G240(1) = AND(G359, G383)
G266(1) = AND(G364, G367, G383, G390)
G229(1) = AND(G366, G396)
G245(1) = AND(G352, G396)
G104BF(1) = NOT(G104)
G97BF(1) = NOT(G97)
G373(1) = NOT(I386)
G392(1) = NOT(I390)
II476(1) = NOT(G384)
I279(1) = NOT(G278)
G249(1) = AND(G366, G66, G397)
G132(1) = NOT(I279)
G374(1) = NOT(G373)
G393(1) = NOT(G392)
G224(1) = NOT(II476)
G282(1) = OR(G233, G249, G263)
G253(1) = AND(G356, G373, G375)
I533(1) = AND(G365, G367, G373)
G227(1) = AND(G366, G392)
G243(1) = AND(G392, G361)
I306(1) = NOT(G282)
G268(1) = OR(G224, G240)
G265(1) = AND(G375, G390, I533)
G236(1) = AND(G374, G376)
G237(1) = AND(G374, G375)
G252(1) = AND(G355, G374, G375)
II527(1) = AND(G366, G64, G393)
G286(1) = OR(G237, G253)
G285(1) = OR(G236, G252)
II208(1) = NOT(G268)
I308(1) = NOT(I306)
I307(1) = NAND(G282, I306)
I334(1) = NOT(G286)
I327(1) = NOT(G285)
I210(1) = NOT(II208)
G136(1) = NAND(I307, I308)
I209(1) = NAND(G268, II208)
G122(1) = NAND(I209, I210)
I336(1) = NOT(I334)
I329(1) = NOT(I327)
I442(1) = NOT(G136)
II335(1) = NAND(G286, I334)
I328(1) = NAND(G285, I327)
G139(1) = NAND(I328, I329)
G140(1) = NAND(II335, I336)
G331(1) = NOT(I442)
G88(1) = AND(G331, G24)
G88BF(1) = NOT(G88)
I414(1) = NOT(G88)
G178(1) = NOT(I414)
I449(1) = NOT(G178)
G179(1) = NOT(I449)
I452(1) = NOT(G179)
G357(1) = NOT(I452)
G358(1) = NOT(G357)
G112(1) = NOT(G358)
G212(1) = NAND(G379, G358)
G335(1) = AND(G112, G113)
G306(1) = AND(G212, G213)
I460(1) = NOT(G335)
I463(1) = NOT(G335)
I466(1) = NOT(G306)
I469(1) = NOT(G306)
G190(1) = NOT(I460)
G336(1) = NOT(I463)
G158(1) = NOT(I466)
G307(1) = NOT(I469)
I472(1) = NOT(G190)
I476(1) = NOT(G158)
G99(1) = AND(G336, G34)
G395(1) = NOT(G158)
G105(1) = AND(G307, G16)
G277(1) = AND(G366, G158, G397)
G228(1) = AND(G366, G158)
G244(1) = AND(G158, G362)
G105BF(1) = NOT(G105)
G99BF(1) = NOT(G99)
G262(1) = AND(G366, G392, G395, G397)
G394(1) = NOT(I476)
G377(1) = NOT(I472)
II272(1) = NOT(G277)
G276(1) = AND(G366, G392, G395, G397)
I515(1) = AND(G393, G395, G397)
G261(1) = AND(G395, G397, II527)
G131(1) = NOT(II272)
G378(1) = NOT(G377)
I265(1) = NOT(G276)
G280(1) = OR(G231, G247, G261)
G251(1) = AND(G358, G377, G381)
I512(1) = AND(G364, G368, G377)
II538(1) = AND(G377, G381, G383, G387)
G130(1) = NOT(I265)
I292(1) = NOT(G280)
G256(1) = AND(G381, G390, I512)
G230(1) = AND(G378, G382)
G235(1) = AND(G378, G381)
G246(1) = AND(G357, G378, G381)
G284(1) = OR(G235, G251)
G279(1) = OR(G230, G246)
I294(1) = NOT(I292)
I293(1) = NAND(G280, I292)
I320(1) = NOT(G284)
I285(1) = NOT(G279)
G134(1) = NAND(I293, I294)
I322(1) = NOT(I320)
II287(1) = NOT(I285)
I517(1) = NOT(G134)
II321(1) = NAND(G284, I320)
I286(1) = NAND(G279, I285)
G133(1) = NAND(I286, II287)
G138(1) = NAND(II321, I322)
G327(1) = NOT(I517)
G86(1) = AND(G327, G22)
G86BF(1) = NOT(G86)
I398(1) = NOT(G86)
G168(1) = NOT(I398)
I524(1) = NOT(G168)
G169(1) = NOT(I524)
I527(1) = NOT(G169)
G353(1) = NOT(I527)
G354(1) = NOT(G353)
G120(1) = NOT(G354)
G208(1) = NAND(G379, G354)
G347(1) = AND(G120, G121)
G300(1) = AND(G208, G209)
I535(1) = NOT(G347)
I538(1) = NOT(G347)
I541(1) = NOT(G300)
I544(1) = NOT(G300)
G206(1) = NOT(I535)
G348(1) = NOT(I538)
G150(1) = NOT(I541)
G301(1) = NOT(I544)
I547(1) = NOT(G206)
I551(1) = NOT(G150)
G95(1) = AND(G348, G30)
G391(1) = NOT(G150)
G103(1) = AND(G301, G14)
G226(1) = AND(G366, G150)
G242(1) = AND(G150, G363)
I553(1) = AND(G366, G150, G393)
G103BF(1) = NOT(G103)
G95BF(1) = NOT(G95)
G380(1) = NOT(I551)
G369(1) = NOT(I547)
G275(1) = AND(G395, G397, I553)
I518(1) = AND(G391, G395, G397)
I521(1) = AND(G391, G393, G397)
II524(1) = AND(G352, G391, G393)
G370(1) = NOT(G369)
I258(1) = NOT(G275)
I495(1) = AND(G365, G368, G369)
G255(1) = AND(G354, G369, G371)
G257(1) = AND(G363, G369, G371, I515)
I537(1) = AND(G369, G371, G373, G375)
G258(1) = AND(G361, G373, G375, I518)
G259(1) = AND(G362, G377, G381, I521)
G260(1) = AND(G395, G383, II524)
G129(1) = NOT(I258)
G271(1) = OR(G226, G242, G257)
G272(1) = OR(G227, G243, G258)
G273(1) = OR(G228, G244, G259)
G274(1) = OR(G229, G245, G260)
G241(1) = AND(G371, G390, I495)
G267(1) = AND(I537, II538)
G238(1) = AND(G370, G372)
G239(1) = AND(G370, G371)
G254(1) = AND(G353, G370, G371)
I230(1) = NOT(G271)
G288(1) = OR(G239, G255)
G287(1) = OR(G238, G254)
I237(1) = NOT(G272)
I244(1) = NOT(G273)
I251(1) = NOT(G274)
I546(1) = OR(G225, G241, G256)
G125(1) = NOT(I230)
G126(1) = NOT(I237)
G127(1) = NOT(I244)
G128(1) = NOT(I251)
I348(1) = NOT(G288)
II341(1) = NOT(G287)
G270(1) = OR(G265, G266, G267, I546)
I222(1) = NOT(G270)
I350(1) = NOT(I348)
I343(1) = NOT(II341)
I349(1) = NAND(G288, I348)
I342(1) = NAND(G287, II341)
G141(1) = NAND(I342, I343)
G142(1) = NAND(I349, I350)
I224(1) = NOT(I222)
I223(1) = NAND(G270, I222)
G124(1) = NAND(I223, I224)
I608(1) = NOT(G124)
G298(1) = NOT(I608)
G90(1) = AND(G298, G26)
