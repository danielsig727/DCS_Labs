# INPUT 36
# OUTPUT 7
# NOT 49
# AND 138
# OR 18
# BUF 40
INPUT(1GAT_0)
INPUT(4GAT_1)
INPUT(8GAT_2)
INPUT(11GAT_3)
INPUT(14GAT_4)
INPUT(17GAT_5)
INPUT(21GAT_6)
INPUT(24GAT_7)
INPUT(27GAT_8)
INPUT(30GAT_9)
INPUT(34GAT_10)
INPUT(37GAT_11)
INPUT(40GAT_12)
INPUT(43GAT_13)
INPUT(47GAT_14)
INPUT(50GAT_15)
INPUT(53GAT_16)
INPUT(56GAT_17)
INPUT(60GAT_18)
INPUT(63GAT_19)
INPUT(66GAT_20)
INPUT(69GAT_21)
INPUT(73GAT_22)
INPUT(76GAT_23)
INPUT(79GAT_24)
INPUT(82GAT_25)
INPUT(86GAT_26)
INPUT(89GAT_27)
INPUT(92GAT_28)
INPUT(95GAT_29)
INPUT(99GAT_30)
INPUT(102GAT_31)
INPUT(105GAT_32)
INPUT(108GAT_33)
INPUT(112GAT_34)
INPUT(115GAT_35)
OUTPUT(223GAT_84)
OUTPUT(329GAT_133)
OUTPUT(370GAT_163)
OUTPUT(421GAT_188)
OUTPUT(430GAT_193)
OUTPUT(431GAT_194)
OUTPUT(432GAT_195)
151GAT_36(1) = BUF(108GAT_33)
150GAT_37(1) = BUF(102GAT_31)
147GAT_38(1) = BUF(95GAT_29)
146GAT_39(1) = BUF(89GAT_27)
143GAT_40(1) = BUF(82GAT_25)
142GAT_41(1) = BUF(76GAT_23)
139GAT_42(1) = BUF(69GAT_21)
138GAT_43(1) = BUF(63GAT_19)
135GAT_44(1) = BUF(56GAT_17)
134GAT_45(1) = BUF(50GAT_15)
131GAT_46(1) = BUF(43GAT_13)
130GAT_47(1) = BUF(37GAT_11)
127GAT_48(1) = BUF(30GAT_9)
126GAT_49(1) = BUF(24GAT_7)
123GAT_50(1) = BUF(17GAT_5)
122GAT_51(1) = BUF(11GAT_3)
119GAT_52(1) = BUF(4GAT_1)
118GAT_53(1) = BUF(1GAT_0)
115GAT_35b(1) = NOT(115GAT_35)
112GAT_34b(1) = NOT(112GAT_34)
105GAT_32b(1) = NOT(105GAT_32)
99GAT_30b(1) = NOT(99GAT_30)
92GAT_28b(1) = NOT(92GAT_28)
86GAT_26b(1) = NOT(86GAT_26)
79GAT_24b(1) = NOT(79GAT_24)
73GAT_22b(1) = NOT(73GAT_22)
66GAT_20b(1) = NOT(66GAT_20)
60GAT_18b(1) = NOT(60GAT_18)
53GAT_16b(1) = NOT(53GAT_16)
47GAT_14b(1) = NOT(47GAT_14)
40GAT_12b(1) = NOT(40GAT_12)
34GAT_10b(1) = NOT(34GAT_10)
27GAT_8b(1) = NOT(27GAT_8)
21GAT_6b(1) = NOT(21GAT_6)
14GAT_4b(1) = NOT(14GAT_4)
8GAT_2b(1) = NOT(8GAT_2)
151GAT_36b(1) = NOT(151GAT_36)
180GAT_56(1) = AND(108GAT_33, 150GAT_37)
147GAT_38b(1) = NOT(147GAT_38)
177GAT_59(1) = AND(95GAT_29, 146GAT_39)
143GAT_40b(1) = NOT(143GAT_40)
174GAT_62(1) = AND(82GAT_25, 142GAT_41)
139GAT_42b(1) = NOT(139GAT_42)
171GAT_65(1) = AND(69GAT_21, 138GAT_43)
135GAT_44b(1) = NOT(135GAT_44)
168GAT_68(1) = AND(56GAT_17, 134GAT_45)
131GAT_46b(1) = NOT(131GAT_46)
165GAT_71(1) = AND(43GAT_13, 130GAT_47)
127GAT_48b(1) = NOT(127GAT_48)
162GAT_74(1) = AND(30GAT_9, 126GAT_49)
123GAT_50b(1) = NOT(123GAT_50)
159GAT_77(1) = AND(17GAT_5, 122GAT_51)
119GAT_52b(1) = NOT(119GAT_52)
154GAT_80(1) = AND(4GAT_1, 118GAT_53)
199GAT_81(1) = AND(180GAT_56, 177GAT_59, 174GAT_62, 171GAT_65, 168GAT_68, 165GAT_71, 162GAT_74, 159GAT_77, 154GAT_80)
198GAT_54(1) = AND(151GAT_36b, 115GAT_35b)
197GAT_55(1) = AND(151GAT_36b, 112GAT_34b)
196GAT_57(1) = AND(147GAT_38b, 105GAT_32b)
195GAT_58(1) = AND(147GAT_38b, 99GAT_30b)
194GAT_60(1) = AND(143GAT_40b, 92GAT_28b)
193GAT_61(1) = AND(143GAT_40b, 86GAT_26b)
192GAT_63(1) = AND(139GAT_42b, 79GAT_24b)
191GAT_64(1) = AND(139GAT_42b, 73GAT_22b)
190GAT_66(1) = AND(135GAT_44b, 66GAT_20b)
189GAT_67(1) = AND(135GAT_44b, 60GAT_18b)
188GAT_69(1) = AND(131GAT_46b, 53GAT_16b)
187GAT_70(1) = AND(131GAT_46b, 47GAT_14b)
186GAT_72(1) = AND(127GAT_48b, 40GAT_12b)
185GAT_73(1) = AND(127GAT_48b, 34GAT_10b)
184GAT_75(1) = AND(123GAT_50b, 27GAT_8b)
183GAT_76(1) = AND(123GAT_50b, 21GAT_6b)
158GAT_78(1) = AND(119GAT_52b, 14GAT_4b)
157GAT_79(1) = AND(119GAT_52b, 8GAT_2b)
180GAT_56b(1) = NOT(180GAT_56)
177GAT_59b(1) = NOT(177GAT_59)
174GAT_62b(1) = NOT(174GAT_62)
171GAT_65b(1) = NOT(171GAT_65)
168GAT_68b(1) = NOT(168GAT_68)
165GAT_71b(1) = NOT(165GAT_71)
162GAT_74b(1) = NOT(162GAT_74)
159GAT_77b(1) = NOT(159GAT_77)
154GAT_80b(1) = NOT(154GAT_80)
223GAT_84(1) = BUF(199GAT_81)
203GAT_82(1) = BUF(199GAT_81)
213GAT_83(1) = BUF(199GAT_81)
internal__52(1) = AND(180GAT_56b, 203GAT_82)
203GAT_82b(1) = NOT(203GAT_82)
259GAT_86(1) = AND(102GAT_31, 213GAT_83)
internal__56(1) = AND(177GAT_59b, 203GAT_82)
258GAT_88(1) = AND(89GAT_27, 213GAT_83)
internal__60(1) = AND(174GAT_62b, 203GAT_82)
257GAT_90(1) = AND(76GAT_23, 213GAT_83)
internal__64(1) = AND(171GAT_65b, 203GAT_82)
256GAT_92(1) = AND(63GAT_19, 213GAT_83)
internal__68(1) = AND(168GAT_68b, 203GAT_82)
255GAT_94(1) = AND(50GAT_15, 213GAT_83)
internal__72(1) = AND(165GAT_71b, 203GAT_82)
254GAT_96(1) = AND(37GAT_11, 213GAT_83)
internal__76(1) = AND(162GAT_74b, 203GAT_82)
250GAT_98(1) = AND(24GAT_7, 213GAT_83)
internal__80(1) = AND(159GAT_77b, 203GAT_82)
246GAT_100(1) = AND(11GAT_3, 213GAT_83)
internal__84(1) = AND(154GAT_80b, 203GAT_82)
242GAT_102(1) = AND(213GAT_83, 1GAT_0)
internal__51(1) = AND(180GAT_56, 203GAT_82b)
internal__55(1) = AND(177GAT_59, 203GAT_82b)
internal__59(1) = AND(174GAT_62, 203GAT_82b)
internal__63(1) = AND(171GAT_65, 203GAT_82b)
internal__67(1) = AND(168GAT_68, 203GAT_82b)
internal__71(1) = AND(165GAT_71, 203GAT_82b)
internal__75(1) = AND(162GAT_74, 203GAT_82b)
internal__79(1) = AND(159GAT_77, 203GAT_82b)
internal__83(1) = AND(154GAT_80, 203GAT_82b)
251GAT_85(1) = OR(internal__52, internal__51)
247GAT_87(1) = OR(internal__56, internal__55)
243GAT_89(1) = OR(internal__60, internal__59)
239GAT_91(1) = OR(internal__64, internal__63)
236GAT_93(1) = OR(internal__68, internal__67)
233GAT_95(1) = OR(internal__72, internal__71)
230GAT_97(1) = OR(internal__76, internal__75)
227GAT_99(1) = OR(internal__80, internal__79)
224GAT_101(1) = OR(internal__84, internal__83)
295GAT_103(1) = AND(198GAT_54, 251GAT_85)
285GAT_104(1) = AND(197GAT_55, 251GAT_85)
294GAT_105(1) = AND(196GAT_57, 247GAT_87)
282GAT_106(1) = AND(195GAT_58, 247GAT_87)
293GAT_107(1) = AND(194GAT_60, 243GAT_89)
279GAT_108(1) = AND(193GAT_61, 243GAT_89)
292GAT_109(1) = AND(192GAT_63, 239GAT_91)
276GAT_110(1) = AND(191GAT_64, 239GAT_91)
291GAT_111(1) = AND(190GAT_66, 236GAT_93)
273GAT_112(1) = AND(189GAT_67, 236GAT_93)
290GAT_113(1) = AND(188GAT_69, 233GAT_95)
270GAT_114(1) = AND(187GAT_70, 233GAT_95)
289GAT_115(1) = AND(186GAT_72, 230GAT_97)
267GAT_116(1) = AND(185GAT_73, 230GAT_97)
288GAT_117(1) = AND(184GAT_75, 227GAT_99)
264GAT_118(1) = AND(183GAT_76, 227GAT_99)
263GAT_119(1) = AND(158GAT_78, 224GAT_101)
260GAT_120(1) = AND(157GAT_79, 224GAT_101)
296GAT_122(1) = AND(285GAT_104, 282GAT_106, 279GAT_108, 276GAT_110, 273GAT_112, 270GAT_114, 267GAT_116, 264GAT_118, 260GAT_120)
308GAT_121(1) = BUF(295GAT_103)
307GAT_123(1) = BUF(294GAT_105)
306GAT_124(1) = BUF(293GAT_107)
305GAT_125(1) = BUF(292GAT_109)
304GAT_126(1) = BUF(291GAT_111)
303GAT_127(1) = BUF(290GAT_113)
302GAT_128(1) = BUF(289GAT_115)
301GAT_129(1) = BUF(288GAT_117)
300GAT_130(1) = BUF(263GAT_119)
285GAT_104b(1) = NOT(285GAT_104)
282GAT_106b(1) = NOT(282GAT_106)
279GAT_108b(1) = NOT(279GAT_108)
276GAT_110b(1) = NOT(276GAT_110)
273GAT_112b(1) = NOT(273GAT_112)
270GAT_114b(1) = NOT(270GAT_114)
267GAT_116b(1) = NOT(267GAT_116)
264GAT_118b(1) = NOT(264GAT_118)
260GAT_120b(1) = NOT(260GAT_120)
329GAT_133(1) = BUF(296GAT_122)
309GAT_131(1) = BUF(296GAT_122)
319GAT_132(1) = BUF(296GAT_122)
347GAT_134(1) = AND(112GAT_34, 319GAT_132)
internal__120(1) = AND(285GAT_104b, 309GAT_131)
309GAT_131b(1) = NOT(309GAT_131)
346GAT_136(1) = AND(99GAT_30, 319GAT_132)
internal__124(1) = AND(282GAT_106b, 309GAT_131)
345GAT_138(1) = AND(86GAT_26, 319GAT_132)
internal__128(1) = AND(279GAT_108b, 309GAT_131)
344GAT_140(1) = AND(73GAT_22, 319GAT_132)
internal__132(1) = AND(276GAT_110b, 309GAT_131)
342GAT_142(1) = AND(60GAT_18, 319GAT_132)
internal__136(1) = AND(273GAT_112b, 309GAT_131)
340GAT_144(1) = AND(47GAT_14, 319GAT_132)
internal__140(1) = AND(270GAT_114b, 309GAT_131)
338GAT_146(1) = AND(34GAT_10, 319GAT_132)
internal__144(1) = AND(267GAT_116b, 309GAT_131)
336GAT_148(1) = AND(21GAT_6, 319GAT_132)
internal__148(1) = AND(264GAT_118b, 309GAT_131)
334GAT_150(1) = AND(319GAT_132, 8GAT_2)
internal__152(1) = AND(260GAT_120b, 309GAT_131)
internal__119(1) = AND(285GAT_104, 309GAT_131b)
internal__123(1) = AND(282GAT_106, 309GAT_131b)
internal__127(1) = AND(279GAT_108, 309GAT_131b)
internal__131(1) = AND(276GAT_110, 309GAT_131b)
internal__135(1) = AND(273GAT_112, 309GAT_131b)
internal__139(1) = AND(270GAT_114, 309GAT_131b)
internal__143(1) = AND(267GAT_116, 309GAT_131b)
internal__147(1) = AND(264GAT_118, 309GAT_131b)
internal__151(1) = AND(260GAT_120, 309GAT_131b)
343GAT_135(1) = OR(internal__120, internal__119)
341GAT_137(1) = OR(internal__124, internal__123)
339GAT_139(1) = OR(internal__128, internal__127)
337GAT_141(1) = OR(internal__132, internal__131)
335GAT_143(1) = OR(internal__136, internal__135)
333GAT_145(1) = OR(internal__140, internal__139)
332GAT_147(1) = OR(internal__144, internal__143)
331GAT_149(1) = OR(internal__148, internal__147)
330GAT_151(1) = OR(internal__152, internal__151)
356GAT_152(1) = AND(308GAT_121, 343GAT_135)
355GAT_153(1) = AND(307GAT_123, 341GAT_137)
354GAT_154(1) = AND(306GAT_124, 339GAT_139)
353GAT_155(1) = AND(305GAT_125, 337GAT_141)
352GAT_156(1) = AND(304GAT_126, 335GAT_143)
351GAT_157(1) = AND(303GAT_127, 333GAT_145)
350GAT_158(1) = AND(302GAT_128, 332GAT_147)
349GAT_159(1) = AND(301GAT_129, 331GAT_149)
348GAT_160(1) = AND(300GAT_130, 330GAT_151)
357GAT_161(1) = AND(356GAT_152, 355GAT_153, 354GAT_154, 353GAT_155, 352GAT_156, 351GAT_157, 350GAT_158, 349GAT_159, 348GAT_160)
370GAT_163(1) = BUF(357GAT_161)
360GAT_162(1) = BUF(357GAT_161)
379GAT_164(1) = AND(115GAT_35, 360GAT_162)
378GAT_165(1) = AND(105GAT_32, 360GAT_162)
377GAT_166(1) = AND(92GAT_28, 360GAT_162)
376GAT_167(1) = AND(79GAT_24, 360GAT_162)
375GAT_168(1) = AND(66GAT_20, 360GAT_162)
374GAT_169(1) = AND(53GAT_16, 360GAT_162)
373GAT_170(1) = AND(40GAT_12, 360GAT_162)
372GAT_171(1) = AND(27GAT_8, 360GAT_162)
371GAT_172(1) = AND(360GAT_162, 14GAT_4)
399GAT_177(1) = AND(56GAT_17, 375GAT_168, 342GAT_142, 255GAT_94)
386GAT_179(1) = AND(30GAT_9, 373GAT_170, 338GAT_146, 250GAT_98)
381GAT_180(1) = AND(17GAT_5, 372GAT_171, 336GAT_148, 246GAT_100)
414GAT_173(1) = AND(108GAT_33, 379GAT_164, 347GAT_134, 259GAT_86)
411GAT_174(1) = AND(95GAT_29, 378GAT_165, 346GAT_136, 258GAT_88)
407GAT_175(1) = AND(82GAT_25, 377GAT_166, 345GAT_138, 257GAT_90)
404GAT_176(1) = AND(69GAT_21, 376GAT_167, 344GAT_140, 256GAT_92)
393GAT_178(1) = AND(43GAT_13, 374GAT_169, 340GAT_144, 254GAT_96)
380GAT_181(1) = AND(371GAT_172, 334GAT_150, 242GAT_102, 4GAT_1)
416GAT_182(1) = AND(414GAT_173, 411GAT_174, 407GAT_175, 404GAT_176, 399GAT_177, 393GAT_178, 386GAT_179, 381GAT_180)
420GAT_183(1) = BUF(411GAT_174)
419GAT_184(1) = BUF(407GAT_175)
418GAT_185(1) = BUF(404GAT_176)
417GAT_186(1) = BUF(393GAT_178)
415GAT_187(1) = BUF(380GAT_181)
416GAT_182b(1) = NOT(416GAT_182)
415GAT_187b(1) = NOT(415GAT_187)
422GAT_192(1) = AND(417GAT_186, 386GAT_179)
428GAT_191(1) = AND(419GAT_184, 393GAT_178, 399GAT_177)
425GAT_190(1) = AND(399GAT_177, 418GAT_185, 393GAT_178, 386GAT_179)
429GAT_189(1) = AND(420GAT_183, 407GAT_175, 393GAT_178, 386GAT_179)
421GAT_188(1) = AND(416GAT_182b, 415GAT_187b)
430GAT_193(1) = AND(399GAT_177, 422GAT_192, 386GAT_179, 381GAT_180)
431GAT_194(1) = AND(428GAT_191, 425GAT_190, 386GAT_179, 381GAT_180)
432GAT_195(1) = AND(429GAT_189, 425GAT_190, 422GAT_192, 381GAT_180)
